`timescale 1ns / 1ps
///////////////////////////////////////////
// ROM table - 2's complement coefficients
// fir_rom2.v: FIR polyphase branch (2)
// 
// Created: 03-Aug-2006 17:33:00
//  from Matlab script fpga_create_rom_verilog.m
//
// J. Shima
//////////////////////////////////////////
module fir_rom2(ADDR, DATA);
    input [8:0] ADDR;
    output signed [15:0] DATA;
    reg signed [15:0] DATA;

    always@(ADDR) begin
        case(ADDR)
          9'b000000000:  DATA = 16'b1111010010101110;    // h1_2=(-0.08844)
          9'b000000001:  DATA = 16'b1111010010011111;    // h2_2=(-0.088898)
          9'b000000010:  DATA = 16'b1111010010010001;    // h3_2=(-0.089325)
          9'b000000011:  DATA = 16'b1111010010000010;    // h4_2=(-0.089783)
          9'b000000100:  DATA = 16'b1111010001110011;    // h5_2=(-0.09024)
          9'b000000101:  DATA = 16'b1111010001100101;    // h6_2=(-0.090668)
          9'b000000110:  DATA = 16'b1111010001010111;    // h7_2=(-0.091095)
          9'b000000111:  DATA = 16'b1111010001001001;    // h8_2=(-0.091522)
          9'b000001000:  DATA = 16'b1111010000111011;    // h9_2=(-0.091949)
          9'b000001001:  DATA = 16'b1111010000101101;    // h10_2=(-0.092377)
          9'b000001010:  DATA = 16'b1111010000011111;    // h11_2=(-0.092804)
          9'b000001011:  DATA = 16'b1111010000010010;    // h12_2=(-0.093201)
          9'b000001100:  DATA = 16'b1111010000000101;    // h13_2=(-0.093597)
          9'b000001101:  DATA = 16'b1111001111111000;    // h14_2=(-0.093994)
          9'b000001110:  DATA = 16'b1111001111101011;    // h15_2=(-0.094391)
          9'b000001111:  DATA = 16'b1111001111011110;    // h16_2=(-0.094788)
          9'b000010000:  DATA = 16'b1111001111010010;    // h17_2=(-0.095154)
          9'b000010001:  DATA = 16'b1111001111000101;    // h18_2=(-0.095551)
          9'b000010010:  DATA = 16'b1111001110111001;    // h19_2=(-0.095917)
          9'b000010011:  DATA = 16'b1111001110101101;    // h20_2=(-0.096283)
          9'b000010100:  DATA = 16'b1111001110100001;    // h21_2=(-0.096649)
          9'b000010101:  DATA = 16'b1111001110010110;    // h22_2=(-0.096985)
          9'b000010110:  DATA = 16'b1111001110001011;    // h23_2=(-0.097321)
          9'b000010111:  DATA = 16'b1111001110000000;    // h24_2=(-0.097656)
          9'b000011000:  DATA = 16'b1111001101110101;    // h25_2=(-0.097992)
          9'b000011001:  DATA = 16'b1111001101101010;    // h26_2=(-0.098328)
          9'b000011010:  DATA = 16'b1111001101011111;    // h27_2=(-0.098663)
          9'b000011011:  DATA = 16'b1111001101010101;    // h28_2=(-0.098969)
          9'b000011100:  DATA = 16'b1111001101001011;    // h29_2=(-0.099274)
          9'b000011101:  DATA = 16'b1111001101000001;    // h30_2=(-0.099579)
          9'b000011110:  DATA = 16'b1111001100111000;    // h31_2=(-0.099854)
          9'b000011111:  DATA = 16'b1111001100101111;    // h32_2=(-0.10013)
          9'b000100000:  DATA = 16'b1111001100100101;    // h33_2=(-0.10043)
          9'b000100001:  DATA = 16'b1111001100011101;    // h34_2=(-0.10068)
          9'b000100010:  DATA = 16'b1111001100010100;    // h35_2=(-0.10095)
          9'b000100011:  DATA = 16'b1111001100001100;    // h36_2=(-0.1012)
          9'b000100100:  DATA = 16'b1111001100000100;    // h37_2=(-0.10144)
          9'b000100101:  DATA = 16'b1111001011111100;    // h38_2=(-0.10168)
          9'b000100110:  DATA = 16'b1111001011110100;    // h39_2=(-0.10193)
          9'b000100111:  DATA = 16'b1111001011101101;    // h40_2=(-0.10214)
          9'b000101000:  DATA = 16'b1111001011100110;    // h41_2=(-0.10236)
          9'b000101001:  DATA = 16'b1111001011011111;    // h42_2=(-0.10257)
          9'b000101010:  DATA = 16'b1111001011011000;    // h43_2=(-0.10278)
          9'b000101011:  DATA = 16'b1111001011010010;    // h44_2=(-0.10297)
          9'b000101100:  DATA = 16'b1111001011001100;    // h45_2=(-0.10315)
          9'b000101101:  DATA = 16'b1111001011000110;    // h46_2=(-0.10333)
          9'b000101110:  DATA = 16'b1111001011000001;    // h47_2=(-0.10349)
          9'b000101111:  DATA = 16'b1111001010111100;    // h48_2=(-0.10364)
          9'b000110000:  DATA = 16'b1111001010110111;    // h49_2=(-0.10379)
          9'b000110001:  DATA = 16'b1111001010110010;    // h50_2=(-0.10394)
          9'b000110010:  DATA = 16'b1111001010101110;    // h51_2=(-0.10406)
          9'b000110011:  DATA = 16'b1111001010101010;    // h52_2=(-0.10419)
          9'b000110100:  DATA = 16'b1111001010100110;    // h53_2=(-0.10431)
          9'b000110101:  DATA = 16'b1111001010100011;    // h54_2=(-0.1044)
          9'b000110110:  DATA = 16'b1111001010100000;    // h55_2=(-0.10449)
          9'b000110111:  DATA = 16'b1111001010011101;    // h56_2=(-0.10458)
          9'b000111000:  DATA = 16'b1111001010011011;    // h57_2=(-0.10464)
          9'b000111001:  DATA = 16'b1111001010011001;    // h58_2=(-0.10471)
          9'b000111010:  DATA = 16'b1111001010010111;    // h59_2=(-0.10477)
          9'b000111011:  DATA = 16'b1111001010010101;    // h60_2=(-0.10483)
          9'b000111100:  DATA = 16'b1111001010010100;    // h61_2=(-0.10486)
          9'b000111101:  DATA = 16'b1111001010010011;    // h62_2=(-0.10489)
          9'b000111110:  DATA = 16'b1111001010010011;    // h63_2=(-0.10489)
          9'b000111111:  DATA = 16'b1111001010010011;    // h64_2=(-0.10489)
          9'b001000000:  DATA = 16'b1111001010010011;    // h65_2=(-0.10489)
          9'b001000001:  DATA = 16'b1111001010010011;    // h66_2=(-0.10489)
          9'b001000010:  DATA = 16'b1111001010010100;    // h67_2=(-0.10486)
          9'b001000011:  DATA = 16'b1111001010010101;    // h68_2=(-0.10483)
          9'b001000100:  DATA = 16'b1111001010010111;    // h69_2=(-0.10477)
          9'b001000101:  DATA = 16'b1111001010011001;    // h70_2=(-0.10471)
          9'b001000110:  DATA = 16'b1111001010011011;    // h71_2=(-0.10464)
          9'b001000111:  DATA = 16'b1111001010011110;    // h72_2=(-0.10455)
          9'b001001000:  DATA = 16'b1111001010100001;    // h73_2=(-0.10446)
          9'b001001001:  DATA = 16'b1111001010100100;    // h74_2=(-0.10437)
          9'b001001010:  DATA = 16'b1111001010101000;    // h75_2=(-0.10425)
          9'b001001011:  DATA = 16'b1111001010101100;    // h76_2=(-0.10413)
          9'b001001100:  DATA = 16'b1111001010110000;    // h77_2=(-0.104)
          9'b001001101:  DATA = 16'b1111001010110101;    // h78_2=(-0.10385)
          9'b001001110:  DATA = 16'b1111001010111010;    // h79_2=(-0.1037)
          9'b001001111:  DATA = 16'b1111001011000000;    // h80_2=(-0.10352)
          9'b001010000:  DATA = 16'b1111001011000110;    // h81_2=(-0.10333)
          9'b001010001:  DATA = 16'b1111001011001100;    // h82_2=(-0.10315)
          9'b001010010:  DATA = 16'b1111001011010011;    // h83_2=(-0.10294)
          9'b001010011:  DATA = 16'b1111001011011010;    // h84_2=(-0.10272)
          9'b001010100:  DATA = 16'b1111001011100010;    // h85_2=(-0.10248)
          9'b001010101:  DATA = 16'b1111001011101010;    // h86_2=(-0.10223)
          9'b001010110:  DATA = 16'b1111001011110010;    // h87_2=(-0.10199)
          9'b001010111:  DATA = 16'b1111001011111011;    // h88_2=(-0.10172)
          9'b001011000:  DATA = 16'b1111001100000100;    // h89_2=(-0.10144)
          9'b001011001:  DATA = 16'b1111001100001110;    // h90_2=(-0.10114)
          9'b001011010:  DATA = 16'b1111001100011000;    // h91_2=(-0.10083)
          9'b001011011:  DATA = 16'b1111001100100010;    // h92_2=(-0.10052)
          9'b001011100:  DATA = 16'b1111001100101101;    // h93_2=(-0.10019)
          9'b001011101:  DATA = 16'b1111001100111000;    // h94_2=(-0.099854)
          9'b001011110:  DATA = 16'b1111001101000100;    // h95_2=(-0.099487)
          9'b001011111:  DATA = 16'b1111001101010000;    // h96_2=(-0.099121)
          9'b001100000:  DATA = 16'b1111001101011101;    // h97_2=(-0.098724)
          9'b001100001:  DATA = 16'b1111001101101010;    // h98_2=(-0.098328)
          9'b001100010:  DATA = 16'b1111001101110111;    // h99_2=(-0.097931)
          9'b001100011:  DATA = 16'b1111001110000101;    // h100_2=(-0.097504)
          9'b001100100:  DATA = 16'b1111001110010011;    // h101_2=(-0.097076)
          9'b001100101:  DATA = 16'b1111001110100010;    // h102_2=(-0.096619)
          9'b001100110:  DATA = 16'b1111001110110001;    // h103_2=(-0.096161)
          9'b001100111:  DATA = 16'b1111001111000001;    // h104_2=(-0.095673)
          9'b001101000:  DATA = 16'b1111001111010001;    // h105_2=(-0.095184)
          9'b001101001:  DATA = 16'b1111001111100010;    // h106_2=(-0.094666)
          9'b001101010:  DATA = 16'b1111001111110011;    // h107_2=(-0.094147)
          9'b001101011:  DATA = 16'b1111010000000100;    // h108_2=(-0.093628)
          9'b001101100:  DATA = 16'b1111010000010110;    // h109_2=(-0.093079)
          9'b001101101:  DATA = 16'b1111010000101000;    // h110_2=(-0.092529)
          9'b001101110:  DATA = 16'b1111010000111011;    // h111_2=(-0.091949)
          9'b001101111:  DATA = 16'b1111010001001111;    // h112_2=(-0.091339)
          9'b001110000:  DATA = 16'b1111010001100010;    // h113_2=(-0.090759)
          9'b001110001:  DATA = 16'b1111010001110111;    // h114_2=(-0.090118)
          9'b001110010:  DATA = 16'b1111010010001100;    // h115_2=(-0.089478)
          9'b001110011:  DATA = 16'b1111010010100001;    // h116_2=(-0.088837)
          9'b001110100:  DATA = 16'b1111010010110111;    // h117_2=(-0.088165)
          9'b001110101:  DATA = 16'b1111010011001101;    // h118_2=(-0.087494)
          9'b001110110:  DATA = 16'b1111010011100011;    // h119_2=(-0.086823)
          9'b001110111:  DATA = 16'b1111010011111011;    // h120_2=(-0.08609)
          9'b001111000:  DATA = 16'b1111010100010010;    // h121_2=(-0.085388)
          9'b001111001:  DATA = 16'b1111010100101011;    // h122_2=(-0.084625)
          9'b001111010:  DATA = 16'b1111010101000011;    // h123_2=(-0.083893)
          9'b001111011:  DATA = 16'b1111010101011100;    // h124_2=(-0.08313)
          9'b001111100:  DATA = 16'b1111010101110110;    // h125_2=(-0.082336)
          9'b001111101:  DATA = 16'b1111010110010000;    // h126_2=(-0.081543)
          9'b001111110:  DATA = 16'b1111010110101011;    // h127_2=(-0.080719)
          9'b001111111:  DATA = 16'b1111010111000110;    // h128_2=(-0.079895)
          9'b010000000:  DATA = 16'b1111010111100010;    // h129_2=(-0.079041)
          9'b010000001:  DATA = 16'b1111010111111110;    // h130_2=(-0.078186)
          9'b010000010:  DATA = 16'b1111011000011011;    // h131_2=(-0.077301)
          9'b010000011:  DATA = 16'b1111011000111000;    // h132_2=(-0.076416)
          9'b010000100:  DATA = 16'b1111011001010110;    // h133_2=(-0.0755)
          9'b010000101:  DATA = 16'b1111011001110100;    // h134_2=(-0.074585)
          9'b010000110:  DATA = 16'b1111011010010011;    // h135_2=(-0.073639)
          9'b010000111:  DATA = 16'b1111011010110010;    // h136_2=(-0.072693)
          9'b010001000:  DATA = 16'b1111011011010010;    // h137_2=(-0.071716)
          9'b010001001:  DATA = 16'b1111011011110010;    // h138_2=(-0.07074)
          9'b010001010:  DATA = 16'b1111011100010011;    // h139_2=(-0.069733)
          9'b010001011:  DATA = 16'b1111011100110101;    // h140_2=(-0.068695)
          9'b010001100:  DATA = 16'b1111011101010111;    // h141_2=(-0.067657)
          9'b010001101:  DATA = 16'b1111011101111001;    // h142_2=(-0.06662)
          9'b010001110:  DATA = 16'b1111011110011100;    // h143_2=(-0.065552)
          9'b010001111:  DATA = 16'b1111011111000000;    // h144_2=(-0.064453)
          9'b010010000:  DATA = 16'b1111011111100100;    // h145_2=(-0.063354)
          9'b010010001:  DATA = 16'b1111100000001000;    // h146_2=(-0.062256)
          9'b010010010:  DATA = 16'b1111100000101101;    // h147_2=(-0.061127)
          9'b010010011:  DATA = 16'b1111100001010011;    // h148_2=(-0.059967)
          9'b010010100:  DATA = 16'b1111100001111001;    // h149_2=(-0.058807)
          9'b010010101:  DATA = 16'b1111100010100000;    // h150_2=(-0.057617)
          9'b010010110:  DATA = 16'b1111100011001000;    // h151_2=(-0.056396)
          9'b010010111:  DATA = 16'b1111100011101111;    // h152_2=(-0.055206)
          9'b010011000:  DATA = 16'b1111100100011000;    // h153_2=(-0.053955)
          9'b010011001:  DATA = 16'b1111100101000001;    // h154_2=(-0.052704)
          9'b010011010:  DATA = 16'b1111100101101010;    // h155_2=(-0.051453)
          9'b010011011:  DATA = 16'b1111100110010100;    // h156_2=(-0.050171)
          9'b010011100:  DATA = 16'b1111100110111111;    // h157_2=(-0.048859)
          9'b010011101:  DATA = 16'b1111100111101010;    // h158_2=(-0.047546)
          9'b010011110:  DATA = 16'b1111101000010110;    // h159_2=(-0.046204)
          9'b010011111:  DATA = 16'b1111101001000010;    // h160_2=(-0.044861)
          9'b010100000:  DATA = 16'b1111101001101111;    // h161_2=(-0.043488)
          9'b010100001:  DATA = 16'b1111101010011101;    // h162_2=(-0.042084)
          9'b010100010:  DATA = 16'b1111101011001011;    // h163_2=(-0.04068)
          9'b010100011:  DATA = 16'b1111101011111001;    // h164_2=(-0.039276)
          9'b010100100:  DATA = 16'b1111101100101000;    // h165_2=(-0.037842)
          9'b010100101:  DATA = 16'b1111101101011000;    // h166_2=(-0.036377)
          9'b010100110:  DATA = 16'b1111101110001000;    // h167_2=(-0.034912)
          9'b010100111:  DATA = 16'b1111101110111001;    // h168_2=(-0.033417)
          9'b010101000:  DATA = 16'b1111101111101010;    // h169_2=(-0.031921)
          9'b010101001:  DATA = 16'b1111110000011100;    // h170_2=(-0.030396)
          9'b010101010:  DATA = 16'b1111110001001111;    // h171_2=(-0.028839)
          9'b010101011:  DATA = 16'b1111110010000010;    // h172_2=(-0.027283)
          9'b010101100:  DATA = 16'b1111110010110101;    // h173_2=(-0.025726)
          9'b010101101:  DATA = 16'b1111110011101010;    // h174_2=(-0.024109)
          9'b010101110:  DATA = 16'b1111110100011110;    // h175_2=(-0.022522)
          9'b010101111:  DATA = 16'b1111110101010100;    // h176_2=(-0.020874)
          9'b010110000:  DATA = 16'b1111110110001010;    // h177_2=(-0.019226)
          9'b010110001:  DATA = 16'b1111110111000000;    // h178_2=(-0.017578)
          9'b010110010:  DATA = 16'b1111110111110111;    // h179_2=(-0.0159)
          9'b010110011:  DATA = 16'b1111111000101111;    // h180_2=(-0.014191)
          9'b010110100:  DATA = 16'b1111111001100111;    // h181_2=(-0.012482)
          9'b010110101:  DATA = 16'b1111111010100000;    // h182_2=(-0.010742)
          9'b010110110:  DATA = 16'b1111111011011001;    // h183_2=(-0.0090027)
          9'b010110111:  DATA = 16'b1111111100010011;    // h184_2=(-0.0072327)
          9'b010111000:  DATA = 16'b1111111101001101;    // h185_2=(-0.0054626)
          9'b010111001:  DATA = 16'b1111111110001000;    // h186_2=(-0.0036621)
          9'b010111010:  DATA = 16'b1111111111000100;    // h187_2=(-0.0018311)
          9'b010111011:  DATA = 16'b0000000000000000;    // h188_2=(0)
          9'b010111100:  DATA = 16'b0000000000111101;    // h189_2=(0.0018616)
          9'b010111101:  DATA = 16'b0000000001111010;    // h190_2=(0.0037231)
          9'b010111110:  DATA = 16'b0000000010111000;    // h191_2=(0.0056152)
          9'b010111111:  DATA = 16'b0000000011110110;    // h192_2=(0.0075073)
          9'b011000000:  DATA = 16'b0000000100110101;    // h193_2=(0.0094299)
          9'b011000001:  DATA = 16'b0000000101110101;    // h194_2=(0.011383)
          9'b011000010:  DATA = 16'b0000000110110101;    // h195_2=(0.013336)
          9'b011000011:  DATA = 16'b0000000111110110;    // h196_2=(0.01532)
          9'b011000100:  DATA = 16'b0000001000110111;    // h197_2=(0.017303)
          9'b011000101:  DATA = 16'b0000001001111001;    // h198_2=(0.019318)
          9'b011000110:  DATA = 16'b0000001010111100;    // h199_2=(0.021362)
          9'b011000111:  DATA = 16'b0000001011111111;    // h200_2=(0.023407)
          9'b011001000:  DATA = 16'b0000001101000010;    // h201_2=(0.025452)
          9'b011001001:  DATA = 16'b0000001110000110;    // h202_2=(0.027527)
          9'b011001010:  DATA = 16'b0000001111001011;    // h203_2=(0.029633)
          9'b011001011:  DATA = 16'b0000010000010000;    // h204_2=(0.031738)
          9'b011001100:  DATA = 16'b0000010001010110;    // h205_2=(0.033875)
          9'b011001101:  DATA = 16'b0000010010011100;    // h206_2=(0.036011)
          9'b011001110:  DATA = 16'b0000010011100011;    // h207_2=(0.038177)
          9'b011001111:  DATA = 16'b0000010100101011;    // h208_2=(0.040375)
          9'b011010000:  DATA = 16'b0000010101110011;    // h209_2=(0.042572)
          9'b011010001:  DATA = 16'b0000010110111100;    // h210_2=(0.0448)
          9'b011010010:  DATA = 16'b0000011000000101;    // h211_2=(0.047028)
          9'b011010011:  DATA = 16'b0000011001001111;    // h212_2=(0.049286)
          9'b011010100:  DATA = 16'b0000011010011001;    // h213_2=(0.051544)
          9'b011010101:  DATA = 16'b0000011011100100;    // h214_2=(0.053833)
          9'b011010110:  DATA = 16'b0000011100101111;    // h215_2=(0.056122)
          9'b011010111:  DATA = 16'b0000011101111011;    // h216_2=(0.058441)
          9'b011011000:  DATA = 16'b0000011111001000;    // h217_2=(0.060791)
          9'b011011001:  DATA = 16'b0000100000010101;    // h218_2=(0.063141)
          9'b011011010:  DATA = 16'b0000100001100011;    // h219_2=(0.065521)
          9'b011011011:  DATA = 16'b0000100010110001;    // h220_2=(0.067902)
          9'b011011100:  DATA = 16'b0000100100000000;    // h221_2=(0.070313)
          9'b011011101:  DATA = 16'b0000100101001111;    // h222_2=(0.072723)
          9'b011011110:  DATA = 16'b0000100110011111;    // h223_2=(0.075165)
          9'b011011111:  DATA = 16'b0000100111101111;    // h224_2=(0.077606)
          9'b011100000:  DATA = 16'b0000101001000000;    // h225_2=(0.080078)
          9'b011100001:  DATA = 16'b0000101010010001;    // h226_2=(0.08255)
          9'b011100010:  DATA = 16'b0000101011100011;    // h227_2=(0.085052)
          9'b011100011:  DATA = 16'b0000101100110110;    // h228_2=(0.087585)
          9'b011100100:  DATA = 16'b0000101110001001;    // h229_2=(0.090118)
          9'b011100101:  DATA = 16'b0000101111011101;    // h230_2=(0.092682)
          9'b011100110:  DATA = 16'b0000110000110001;    // h231_2=(0.095245)
          9'b011100111:  DATA = 16'b0000110010000101;    // h232_2=(0.097809)
          9'b011101000:  DATA = 16'b0000110011011011;    // h233_2=(0.10043)
          9'b011101001:  DATA = 16'b0000110100110000;    // h234_2=(0.10303)
          9'b011101010:  DATA = 16'b0000110110000110;    // h235_2=(0.10565)
          9'b011101011:  DATA = 16'b0000110111011101;    // h236_2=(0.10831)
          9'b011101100:  DATA = 16'b0000111000110101;    // h237_2=(0.11099)
          9'b011101101:  DATA = 16'b0000111010001100;    // h238_2=(0.11365)
          9'b011101110:  DATA = 16'b0000111011100101;    // h239_2=(0.11636)
          9'b011101111:  DATA = 16'b0000111100111101;    // h240_2=(0.11905)
          9'b011110000:  DATA = 16'b0000111110010111;    // h241_2=(0.1218)
          9'b011110001:  DATA = 16'b0000111111110001;    // h242_2=(0.12454)
          9'b011110010:  DATA = 16'b0001000001001011;    // h243_2=(0.12729)
          9'b011110011:  DATA = 16'b0001000010100110;    // h244_2=(0.13007)
          9'b011110100:  DATA = 16'b0001000100000001;    // h245_2=(0.13284)
          9'b011110101:  DATA = 16'b0001000101011101;    // h246_2=(0.13565)
          9'b011110110:  DATA = 16'b0001000110111001;    // h247_2=(0.13846)
          9'b011110111:  DATA = 16'b0001001000010110;    // h248_2=(0.1413)
          9'b011111000:  DATA = 16'b0001001001110011;    // h249_2=(0.14413)
          9'b011111001:  DATA = 16'b0001001011010001;    // h250_2=(0.147)
          9'b011111010:  DATA = 16'b0001001100110000;    // h251_2=(0.1499)
          9'b011111011:  DATA = 16'b0001001110001110;    // h252_2=(0.15277)
          9'b011111100:  DATA = 16'b0001001111101110;    // h253_2=(0.1557)
          9'b011111101:  DATA = 16'b0001010001001101;    // h254_2=(0.1586)
          9'b011111110:  DATA = 16'b0001010010101101;    // h255_2=(0.16153)
          9'b011111111:  DATA = 16'b0001010100001110;    // h256_2=(0.16449)
          9'b100000000:  DATA = 16'b0001010101101111;    // h257_2=(0.16745)
          9'b100000001:  DATA = 16'b0001010111010001;    // h258_2=(0.17044)
          9'b100000010:  DATA = 16'b0001011000110011;    // h259_2=(0.17343)
          9'b100000011:  DATA = 16'b0001011010010101;    // h260_2=(0.17642)
          9'b100000100:  DATA = 16'b0001011011111000;    // h261_2=(0.17944)
          9'b100000101:  DATA = 16'b0001011101011100;    // h262_2=(0.1825)
          9'b100000110:  DATA = 16'b0001011111000000;    // h263_2=(0.18555)
          9'b100000111:  DATA = 16'b0001100000100100;    // h264_2=(0.1886)
          9'b100001000:  DATA = 16'b0001100010001001;    // h265_2=(0.19168)
          9'b100001001:  DATA = 16'b0001100011101110;    // h266_2=(0.19476)
          9'b100001010:  DATA = 16'b0001100101010100;    // h267_2=(0.19788)
          9'b100001011:  DATA = 16'b0001100110111010;    // h268_2=(0.20099)
          9'b100001100:  DATA = 16'b0001101000100000;    // h269_2=(0.2041)
          9'b100001101:  DATA = 16'b0001101010000111;    // h270_2=(0.20724)
          9'b100001110:  DATA = 16'b0001101011101110;    // h271_2=(0.21039)
          9'b100001111:  DATA = 16'b0001101101010110;    // h272_2=(0.21356)
          9'b100010000:  DATA = 16'b0001101110111110;    // h273_2=(0.21674)
          9'b100010001:  DATA = 16'b0001110000100111;    // h274_2=(0.21994)
          9'b100010010:  DATA = 16'b0001110010010000;    // h275_2=(0.22314)
          9'b100010011:  DATA = 16'b0001110011111001;    // h276_2=(0.22635)
          9'b100010100:  DATA = 16'b0001110101100011;    // h277_2=(0.22958)
          9'b100010101:  DATA = 16'b0001110111001101;    // h278_2=(0.23282)
          9'b100010110:  DATA = 16'b0001111000111000;    // h279_2=(0.23608)
          9'b100010111:  DATA = 16'b0001111010100011;    // h280_2=(0.23935)
          9'b100011000:  DATA = 16'b0001111100001110;    // h281_2=(0.24261)
          9'b100011001:  DATA = 16'b0001111101111010;    // h282_2=(0.24591)
          9'b100011010:  DATA = 16'b0001111111100110;    // h283_2=(0.24921)
          9'b100011011:  DATA = 16'b0010000001010010;    // h284_2=(0.2525)
          9'b100011100:  DATA = 16'b0010000010111111;    // h285_2=(0.25583)
          9'b100011101:  DATA = 16'b0010000100101100;    // h286_2=(0.25916)
          9'b100011110:  DATA = 16'b0010000110011010;    // h287_2=(0.26251)
          9'b100011111:  DATA = 16'b0010001000001000;    // h288_2=(0.26587)
          9'b100100000:  DATA = 16'b0010001001110110;    // h289_2=(0.26923)
          9'b100100001:  DATA = 16'b0010001011100100;    // h290_2=(0.27258)
          9'b100100010:  DATA = 16'b0010001101010011;    // h291_2=(0.27597)
          9'b100100011:  DATA = 16'b0010001111000011;    // h292_2=(0.27939)
          9'b100100100:  DATA = 16'b0010010000110010;    // h293_2=(0.28278)
          9'b100100101:  DATA = 16'b0010010010100010;    // h294_2=(0.28619)
          9'b100100110:  DATA = 16'b0010010100010010;    // h295_2=(0.28961)
          9'b100100111:  DATA = 16'b0010010110000011;    // h296_2=(0.29306)
          9'b100101000:  DATA = 16'b0010010111110100;    // h297_2=(0.29651)
          9'b100101001:  DATA = 16'b0010011001100101;    // h298_2=(0.29996)
          9'b100101010:  DATA = 16'b0010011011010111;    // h299_2=(0.30344)
          9'b100101011:  DATA = 16'b0010011101001000;    // h300_2=(0.30688)
          9'b100101100:  DATA = 16'b0010011110111010;    // h301_2=(0.31036)
          9'b100101101:  DATA = 16'b0010100000101101;    // h302_2=(0.31387)
          9'b100101110:  DATA = 16'b0010100010011111;    // h303_2=(0.31735)
          9'b100101111:  DATA = 16'b0010100100010010;    // h304_2=(0.32086)
          9'b100110000:  DATA = 16'b0010100110000110;    // h305_2=(0.3244)
          9'b100110001:  DATA = 16'b0010100111111001;    // h306_2=(0.32791)
          9'b100110010:  DATA = 16'b0010101001101101;    // h307_2=(0.33145)
          9'b100110011:  DATA = 16'b0010101011100001;    // h308_2=(0.33499)
          9'b100110100:  DATA = 16'b0010101101010101;    // h309_2=(0.33853)
          9'b100110101:  DATA = 16'b0010101111001010;    // h310_2=(0.3421)
          9'b100110110:  DATA = 16'b0010110000111110;    // h311_2=(0.34564)
          9'b100110111:  DATA = 16'b0010110010110011;    // h312_2=(0.34921)
          9'b100111000:  DATA = 16'b0010110100101000;    // h313_2=(0.35278)
          9'b100111001:  DATA = 16'b0010110110011110;    // h314_2=(0.35638)
          9'b100111010:  DATA = 16'b0010111000010100;    // h315_2=(0.35999)
          9'b100111011:  DATA = 16'b0010111010001010;    // h316_2=(0.36359)
          9'b100111100:  DATA = 16'b0010111100000000;    // h317_2=(0.36719)
          9'b100111101:  DATA = 16'b0010111101110110;    // h318_2=(0.37079)
          9'b100111110:  DATA = 16'b0010111111101100;    // h319_2=(0.37439)
          9'b100111111:  DATA = 16'b0011000001100011;    // h320_2=(0.37802)
          9'b101000000:  DATA = 16'b0011000011011010;    // h321_2=(0.38165)
          9'b101000001:  DATA = 16'b0011000101010001;    // h322_2=(0.38528)
          9'b101000010:  DATA = 16'b0011000111001000;    // h323_2=(0.38892)
          9'b101000011:  DATA = 16'b0011001001000000;    // h324_2=(0.39258)
          9'b101000100:  DATA = 16'b0011001010111000;    // h325_2=(0.39624)
          9'b101000101:  DATA = 16'b0011001100101111;    // h326_2=(0.39987)
          9'b101000110:  DATA = 16'b0011001110100111;    // h327_2=(0.40353)
          9'b101000111:  DATA = 16'b0011010000011111;    // h328_2=(0.4072)
          9'b101001000:  DATA = 16'b0011010010011000;    // h329_2=(0.41089)
          9'b101001001:  DATA = 16'b0011010100010000;    // h330_2=(0.41455)
          9'b101001010:  DATA = 16'b0011010110001001;    // h331_2=(0.41824)
          9'b101001011:  DATA = 16'b0011011000000001;    // h332_2=(0.42191)
          9'b101001100:  DATA = 16'b0011011001111010;    // h333_2=(0.4256)
          9'b101001101:  DATA = 16'b0011011011110011;    // h334_2=(0.42929)
          9'b101001110:  DATA = 16'b0011011101101100;    // h335_2=(0.43298)
          9'b101001111:  DATA = 16'b0011011111100101;    // h336_2=(0.43668)
          9'b101010000:  DATA = 16'b0011100001011110;    // h337_2=(0.44037)
          9'b101010001:  DATA = 16'b0011100011011000;    // h338_2=(0.44409)
          9'b101010010:  DATA = 16'b0011100101010001;    // h339_2=(0.44778)
          9'b101010011:  DATA = 16'b0011100111001011;    // h340_2=(0.45151)
          9'b101010100:  DATA = 16'b0011101001000100;    // h341_2=(0.4552)
          9'b101010101:  DATA = 16'b0011101010111110;    // h342_2=(0.45892)
          9'b101010110:  DATA = 16'b0011101100111000;    // h343_2=(0.46265)
          9'b101010111:  DATA = 16'b0011101110110001;    // h344_2=(0.46634)
          9'b101011000:  DATA = 16'b0011110000101011;    // h345_2=(0.47006)
          9'b101011001:  DATA = 16'b0011110010100101;    // h346_2=(0.47379)
          9'b101011010:  DATA = 16'b0011110100011111;    // h347_2=(0.47751)
          9'b101011011:  DATA = 16'b0011110110011001;    // h348_2=(0.48123)
          9'b101011100:  DATA = 16'b0011111000010011;    // h349_2=(0.48495)
          9'b101011101:  DATA = 16'b0011111010001101;    // h350_2=(0.48868)
          9'b101011110:  DATA = 16'b0011111100000111;    // h351_2=(0.4924)
          9'b101011111:  DATA = 16'b0011111110000001;    // h352_2=(0.49612)
          9'b101100000:  DATA = 16'b0011111111111011;    // h353_2=(0.49985)
          9'b101100001:  DATA = 16'b0100000001110101;    // h354_2=(0.50357)
          9'b101100010:  DATA = 16'b0100000011101111;    // h355_2=(0.50729)
          9'b101100011:  DATA = 16'b0100000101101001;    // h356_2=(0.51102)
          9'b101100100:  DATA = 16'b0100000111100011;    // h357_2=(0.51474)
          9'b101100101:  DATA = 16'b0100001001011101;    // h358_2=(0.51846)
          9'b101100110:  DATA = 16'b0100001011010111;    // h359_2=(0.52219)
          9'b101100111:  DATA = 16'b0100001101010001;    // h360_2=(0.52591)
          9'b101101000:  DATA = 16'b0100001111001011;    // h361_2=(0.52963)
          9'b101101001:  DATA = 16'b0100010001000101;    // h362_2=(0.53336)
          9'b101101010:  DATA = 16'b0100010010111111;    // h363_2=(0.53708)
          9'b101101011:  DATA = 16'b0100010100111001;    // h364_2=(0.5408)
          9'b101101100:  DATA = 16'b0100010110110010;    // h365_2=(0.54449)
          9'b101101101:  DATA = 16'b0100011000101100;    // h366_2=(0.54822)
          9'b101101110:  DATA = 16'b0100011010100101;    // h367_2=(0.55191)
          9'b101101111:  DATA = 16'b0100011100011111;    // h368_2=(0.55563)
          9'b101110000:  DATA = 16'b0100011110011000;    // h369_2=(0.55933)
          9'b101110001:  DATA = 16'b0100100000010001;    // h370_2=(0.56302)
          9'b101110010:  DATA = 16'b0100100010001010;    // h371_2=(0.56671)
          9'b101110011:  DATA = 16'b0100100100000100;    // h372_2=(0.57043)
          9'b101110100:  DATA = 16'b0100100101111100;    // h373_2=(0.5741)
          9'b101110101:  DATA = 16'b0100100111110101;    // h374_2=(0.57779)
          9'b101110110:  DATA = 16'b0100101001101110;    // h375_2=(0.58148)
          default : DATA = 16'b0000000000000000;
        endcase
    end
endmodule

