`timescale 1ns / 1ps
///////////////////////////////////////////
// ROM table - 2's complement coefficients
// fir_rom5.v: FIR polyphase branch (5)
// 
// Created: 03-Aug-2006 17:33:01
//  from Matlab script fpga_create_rom_verilog.m
//
// J. Shima
//////////////////////////////////////////
module fir_rom5(ADDR, DATA);
    input [8:0] ADDR;
    output signed [15:0] DATA;
    reg signed [15:0] DATA;

    always@(ADDR) begin
        case(ADDR)
          9'b000000000:  DATA = 16'b1111010010111101;    // h1_5=(-0.087982)
          9'b000000001:  DATA = 16'b1111010011001101;    // h2_5=(-0.087494)
          9'b000000010:  DATA = 16'b1111010011011100;    // h3_5=(-0.087036)
          9'b000000011:  DATA = 16'b1111010011101100;    // h4_5=(-0.086548)
          9'b000000100:  DATA = 16'b1111010011111011;    // h5_5=(-0.08609)
          9'b000000101:  DATA = 16'b1111010100001011;    // h6_5=(-0.085602)
          9'b000000110:  DATA = 16'b1111010100011011;    // h7_5=(-0.085114)
          9'b000000111:  DATA = 16'b1111010100101011;    // h8_5=(-0.084625)
          9'b000001000:  DATA = 16'b1111010100111011;    // h9_5=(-0.084137)
          9'b000001001:  DATA = 16'b1111010101001100;    // h10_5=(-0.083618)
          9'b000001010:  DATA = 16'b1111010101011100;    // h11_5=(-0.08313)
          9'b000001011:  DATA = 16'b1111010101101100;    // h12_5=(-0.082642)
          9'b000001100:  DATA = 16'b1111010101111101;    // h13_5=(-0.082123)
          9'b000001101:  DATA = 16'b1111010110001110;    // h14_5=(-0.081604)
          9'b000001110:  DATA = 16'b1111010110011111;    // h15_5=(-0.081085)
          9'b000001111:  DATA = 16'b1111010110110000;    // h16_5=(-0.080566)
          9'b000010000:  DATA = 16'b1111010111000001;    // h17_5=(-0.080048)
          9'b000010001:  DATA = 16'b1111010111010010;    // h18_5=(-0.079529)
          9'b000010010:  DATA = 16'b1111010111100011;    // h19_5=(-0.07901)
          9'b000010011:  DATA = 16'b1111010111110100;    // h20_5=(-0.078491)
          9'b000010100:  DATA = 16'b1111011000000110;    // h21_5=(-0.077942)
          9'b000010101:  DATA = 16'b1111011000010111;    // h22_5=(-0.077423)
          9'b000010110:  DATA = 16'b1111011000101000;    // h23_5=(-0.076904)
          9'b000010111:  DATA = 16'b1111011000111010;    // h24_5=(-0.076355)
          9'b000011000:  DATA = 16'b1111011001001100;    // h25_5=(-0.075806)
          9'b000011001:  DATA = 16'b1111011001011110;    // h26_5=(-0.075256)
          9'b000011010:  DATA = 16'b1111011001101111;    // h27_5=(-0.074738)
          9'b000011011:  DATA = 16'b1111011010000001;    // h28_5=(-0.074188)
          9'b000011100:  DATA = 16'b1111011010010011;    // h29_5=(-0.073639)
          9'b000011101:  DATA = 16'b1111011010100101;    // h30_5=(-0.07309)
          9'b000011110:  DATA = 16'b1111011010110111;    // h31_5=(-0.07254)
          9'b000011111:  DATA = 16'b1111011011001001;    // h32_5=(-0.071991)
          9'b000100000:  DATA = 16'b1111011011011100;    // h33_5=(-0.071411)
          9'b000100001:  DATA = 16'b1111011011101110;    // h34_5=(-0.070862)
          9'b000100010:  DATA = 16'b1111011100000000;    // h35_5=(-0.070313)
          9'b000100011:  DATA = 16'b1111011100010011;    // h36_5=(-0.069733)
          9'b000100100:  DATA = 16'b1111011100100101;    // h37_5=(-0.069183)
          9'b000100101:  DATA = 16'b1111011100110111;    // h38_5=(-0.068634)
          9'b000100110:  DATA = 16'b1111011101001010;    // h39_5=(-0.068054)
          9'b000100111:  DATA = 16'b1111011101011100;    // h40_5=(-0.067505)
          9'b000101000:  DATA = 16'b1111011101101111;    // h41_5=(-0.066925)
          9'b000101001:  DATA = 16'b1111011110000001;    // h42_5=(-0.066376)
          9'b000101010:  DATA = 16'b1111011110010100;    // h43_5=(-0.065796)
          9'b000101011:  DATA = 16'b1111011110100111;    // h44_5=(-0.065216)
          9'b000101100:  DATA = 16'b1111011110111001;    // h45_5=(-0.064667)
          9'b000101101:  DATA = 16'b1111011111001100;    // h46_5=(-0.064087)
          9'b000101110:  DATA = 16'b1111011111011111;    // h47_5=(-0.063507)
          9'b000101111:  DATA = 16'b1111011111110001;    // h48_5=(-0.062958)
          9'b000110000:  DATA = 16'b1111100000000100;    // h49_5=(-0.062378)
          9'b000110001:  DATA = 16'b1111100000010111;    // h50_5=(-0.061798)
          9'b000110010:  DATA = 16'b1111100000101010;    // h51_5=(-0.061218)
          9'b000110011:  DATA = 16'b1111100000111100;    // h52_5=(-0.060669)
          9'b000110100:  DATA = 16'b1111100001001111;    // h53_5=(-0.060089)
          9'b000110101:  DATA = 16'b1111100001100010;    // h54_5=(-0.059509)
          9'b000110110:  DATA = 16'b1111100001110101;    // h55_5=(-0.058929)
          9'b000110111:  DATA = 16'b1111100010000111;    // h56_5=(-0.05838)
          9'b000111000:  DATA = 16'b1111100010011010;    // h57_5=(-0.0578)
          9'b000111001:  DATA = 16'b1111100010101101;    // h58_5=(-0.05722)
          9'b000111010:  DATA = 16'b1111100011000000;    // h59_5=(-0.056641)
          9'b000111011:  DATA = 16'b1111100011010010;    // h60_5=(-0.056091)
          9'b000111100:  DATA = 16'b1111100011100101;    // h61_5=(-0.055511)
          9'b000111101:  DATA = 16'b1111100011111000;    // h62_5=(-0.054932)
          9'b000111110:  DATA = 16'b1111100100001011;    // h63_5=(-0.054352)
          9'b000111111:  DATA = 16'b1111100100011101;    // h64_5=(-0.053802)
          9'b001000000:  DATA = 16'b1111100100110000;    // h65_5=(-0.053223)
          9'b001000001:  DATA = 16'b1111100101000011;    // h66_5=(-0.052643)
          9'b001000010:  DATA = 16'b1111100101010101;    // h67_5=(-0.052094)
          9'b001000011:  DATA = 16'b1111100101101000;    // h68_5=(-0.051514)
          9'b001000100:  DATA = 16'b1111100101111011;    // h69_5=(-0.050934)
          9'b001000101:  DATA = 16'b1111100110001101;    // h70_5=(-0.050385)
          9'b001000110:  DATA = 16'b1111100110100000;    // h71_5=(-0.049805)
          9'b001000111:  DATA = 16'b1111100110110010;    // h72_5=(-0.049255)
          9'b001001000:  DATA = 16'b1111100111000101;    // h73_5=(-0.048676)
          9'b001001001:  DATA = 16'b1111100111010111;    // h74_5=(-0.048126)
          9'b001001010:  DATA = 16'b1111100111101010;    // h75_5=(-0.047546)
          9'b001001011:  DATA = 16'b1111100111111100;    // h76_5=(-0.046997)
          9'b001001100:  DATA = 16'b1111101000001110;    // h77_5=(-0.046448)
          9'b001001101:  DATA = 16'b1111101000100001;    // h78_5=(-0.045868)
          9'b001001110:  DATA = 16'b1111101000110011;    // h79_5=(-0.045319)
          9'b001001111:  DATA = 16'b1111101001000101;    // h80_5=(-0.044769)
          9'b001010000:  DATA = 16'b1111101001010111;    // h81_5=(-0.04422)
          9'b001010001:  DATA = 16'b1111101001101001;    // h82_5=(-0.043671)
          9'b001010010:  DATA = 16'b1111101001111011;    // h83_5=(-0.043121)
          9'b001010011:  DATA = 16'b1111101010001101;    // h84_5=(-0.042572)
          9'b001010100:  DATA = 16'b1111101010011111;    // h85_5=(-0.042023)
          9'b001010101:  DATA = 16'b1111101010110001;    // h86_5=(-0.041473)
          9'b001010110:  DATA = 16'b1111101011000011;    // h87_5=(-0.040924)
          9'b001010111:  DATA = 16'b1111101011010101;    // h88_5=(-0.040375)
          9'b001011000:  DATA = 16'b1111101011100111;    // h89_5=(-0.039825)
          9'b001011001:  DATA = 16'b1111101011111000;    // h90_5=(-0.039307)
          9'b001011010:  DATA = 16'b1111101100001010;    // h91_5=(-0.038757)
          9'b001011011:  DATA = 16'b1111101100011100;    // h92_5=(-0.038208)
          9'b001011100:  DATA = 16'b1111101100101101;    // h93_5=(-0.037689)
          9'b001011101:  DATA = 16'b1111101100111110;    // h94_5=(-0.03717)
          9'b001011110:  DATA = 16'b1111101101010000;    // h95_5=(-0.036621)
          9'b001011111:  DATA = 16'b1111101101100001;    // h96_5=(-0.036102)
          9'b001100000:  DATA = 16'b1111101101110010;    // h97_5=(-0.035583)
          9'b001100001:  DATA = 16'b1111101110000100;    // h98_5=(-0.035034)
          9'b001100010:  DATA = 16'b1111101110010101;    // h99_5=(-0.034515)
          9'b001100011:  DATA = 16'b1111101110100110;    // h100_5=(-0.033997)
          9'b001100100:  DATA = 16'b1111101110110111;    // h101_5=(-0.033478)
          9'b001100101:  DATA = 16'b1111101111000111;    // h102_5=(-0.03299)
          9'b001100110:  DATA = 16'b1111101111011000;    // h103_5=(-0.032471)
          9'b001100111:  DATA = 16'b1111101111101001;    // h104_5=(-0.031952)
          9'b001101000:  DATA = 16'b1111101111111010;    // h105_5=(-0.031433)
          9'b001101001:  DATA = 16'b1111110000001010;    // h106_5=(-0.030945)
          9'b001101010:  DATA = 16'b1111110000011011;    // h107_5=(-0.030426)
          9'b001101011:  DATA = 16'b1111110000101011;    // h108_5=(-0.029938)
          9'b001101100:  DATA = 16'b1111110000111011;    // h109_5=(-0.029449)
          9'b001101101:  DATA = 16'b1111110001001011;    // h110_5=(-0.028961)
          9'b001101110:  DATA = 16'b1111110001011100;    // h111_5=(-0.028442)
          9'b001101111:  DATA = 16'b1111110001101100;    // h112_5=(-0.027954)
          9'b001110000:  DATA = 16'b1111110001111100;    // h113_5=(-0.027466)
          9'b001110001:  DATA = 16'b1111110010001011;    // h114_5=(-0.027008)
          9'b001110010:  DATA = 16'b1111110010011011;    // h115_5=(-0.02652)
          9'b001110011:  DATA = 16'b1111110010101011;    // h116_5=(-0.026031)
          9'b001110100:  DATA = 16'b1111110010111010;    // h117_5=(-0.025574)
          9'b001110101:  DATA = 16'b1111110011001010;    // h118_5=(-0.025085)
          9'b001110110:  DATA = 16'b1111110011011001;    // h119_5=(-0.024628)
          9'b001110111:  DATA = 16'b1111110011101001;    // h120_5=(-0.024139)
          9'b001111000:  DATA = 16'b1111110011111000;    // h121_5=(-0.023682)
          9'b001111001:  DATA = 16'b1111110100000111;    // h122_5=(-0.023224)
          9'b001111010:  DATA = 16'b1111110100010110;    // h123_5=(-0.022766)
          9'b001111011:  DATA = 16'b1111110100100101;    // h124_5=(-0.022308)
          9'b001111100:  DATA = 16'b1111110100110100;    // h125_5=(-0.021851)
          9'b001111101:  DATA = 16'b1111110101000010;    // h126_5=(-0.021423)
          9'b001111110:  DATA = 16'b1111110101010001;    // h127_5=(-0.020966)
          9'b001111111:  DATA = 16'b1111110101100000;    // h128_5=(-0.020508)
          9'b010000000:  DATA = 16'b1111110101101110;    // h129_5=(-0.020081)
          9'b010000001:  DATA = 16'b1111110101111100;    // h130_5=(-0.019653)
          9'b010000010:  DATA = 16'b1111110110001011;    // h131_5=(-0.019196)
          9'b010000011:  DATA = 16'b1111110110011001;    // h132_5=(-0.018768)
          9'b010000100:  DATA = 16'b1111110110100111;    // h133_5=(-0.018341)
          9'b010000101:  DATA = 16'b1111110110110101;    // h134_5=(-0.017914)
          9'b010000110:  DATA = 16'b1111110111000010;    // h135_5=(-0.017517)
          9'b010000111:  DATA = 16'b1111110111010000;    // h136_5=(-0.01709)
          9'b010001000:  DATA = 16'b1111110111011110;    // h137_5=(-0.016663)
          9'b010001001:  DATA = 16'b1111110111101011;    // h138_5=(-0.016266)
          9'b010001010:  DATA = 16'b1111110111111001;    // h139_5=(-0.015839)
          9'b010001011:  DATA = 16'b1111111000000110;    // h140_5=(-0.015442)
          9'b010001100:  DATA = 16'b1111111000010011;    // h141_5=(-0.015045)
          9'b010001101:  DATA = 16'b1111111000100000;    // h142_5=(-0.014648)
          9'b010001110:  DATA = 16'b1111111000101101;    // h143_5=(-0.014252)
          9'b010001111:  DATA = 16'b1111111000111010;    // h144_5=(-0.013855)
          9'b010010000:  DATA = 16'b1111111001000111;    // h145_5=(-0.013458)
          9'b010010001:  DATA = 16'b1111111001010011;    // h146_5=(-0.013092)
          9'b010010010:  DATA = 16'b1111111001100000;    // h147_5=(-0.012695)
          9'b010010011:  DATA = 16'b1111111001101100;    // h148_5=(-0.012329)
          9'b010010100:  DATA = 16'b1111111001111001;    // h149_5=(-0.011932)
          9'b010010101:  DATA = 16'b1111111010000101;    // h150_5=(-0.011566)
          9'b010010110:  DATA = 16'b1111111010010001;    // h151_5=(-0.0112)
          9'b010010111:  DATA = 16'b1111111010011101;    // h152_5=(-0.010834)
          9'b010011000:  DATA = 16'b1111111010101001;    // h153_5=(-0.010468)
          9'b010011001:  DATA = 16'b1111111010110100;    // h154_5=(-0.010132)
          9'b010011010:  DATA = 16'b1111111011000000;    // h155_5=(-0.0097656)
          9'b010011011:  DATA = 16'b1111111011001100;    // h156_5=(-0.0093994)
          9'b010011100:  DATA = 16'b1111111011010111;    // h157_5=(-0.0090637)
          9'b010011101:  DATA = 16'b1111111011100010;    // h158_5=(-0.008728)
          9'b010011110:  DATA = 16'b1111111011101101;    // h159_5=(-0.0083923)
          9'b010011111:  DATA = 16'b1111111011111000;    // h160_5=(-0.0080566)
          9'b010100000:  DATA = 16'b1111111100000011;    // h161_5=(-0.0077209)
          9'b010100001:  DATA = 16'b1111111100001110;    // h162_5=(-0.0073853)
          9'b010100010:  DATA = 16'b1111111100011001;    // h163_5=(-0.0070496)
          9'b010100011:  DATA = 16'b1111111100100100;    // h164_5=(-0.0067139)
          9'b010100100:  DATA = 16'b1111111100101110;    // h165_5=(-0.0064087)
          9'b010100101:  DATA = 16'b1111111100111000;    // h166_5=(-0.0061035)
          9'b010100110:  DATA = 16'b1111111101000011;    // h167_5=(-0.0057678)
          9'b010100111:  DATA = 16'b1111111101001101;    // h168_5=(-0.0054626)
          9'b010101000:  DATA = 16'b1111111101010111;    // h169_5=(-0.0051575)
          9'b010101001:  DATA = 16'b1111111101100001;    // h170_5=(-0.0048523)
          9'b010101010:  DATA = 16'b1111111101101011;    // h171_5=(-0.0045471)
          9'b010101011:  DATA = 16'b1111111101110100;    // h172_5=(-0.0042725)
          9'b010101100:  DATA = 16'b1111111101111110;    // h173_5=(-0.0039673)
          9'b010101101:  DATA = 16'b1111111110000111;    // h174_5=(-0.0036926)
          9'b010101110:  DATA = 16'b1111111110010001;    // h175_5=(-0.0033875)
          9'b010101111:  DATA = 16'b1111111110011010;    // h176_5=(-0.0031128)
          9'b010110000:  DATA = 16'b1111111110100011;    // h177_5=(-0.0028381)
          9'b010110001:  DATA = 16'b1111111110101100;    // h178_5=(-0.0025635)
          9'b010110010:  DATA = 16'b1111111110110101;    // h179_5=(-0.0022888)
          9'b010110011:  DATA = 16'b1111111110111110;    // h180_5=(-0.0020142)
          9'b010110100:  DATA = 16'b1111111111000110;    // h181_5=(-0.00177)
          9'b010110101:  DATA = 16'b1111111111001111;    // h182_5=(-0.0014954)
          9'b010110110:  DATA = 16'b1111111111010111;    // h183_5=(-0.0012512)
          9'b010110111:  DATA = 16'b1111111111100000;    // h184_5=(-0.00097656)
          9'b010111000:  DATA = 16'b1111111111101000;    // h185_5=(-0.00073242)
          9'b010111001:  DATA = 16'b1111111111110000;    // h186_5=(-0.00048828)
          9'b010111010:  DATA = 16'b1111111111111000;    // h187_5=(-0.00024414)
          9'b010111011:  DATA = 16'b0000000000000000;    // h188_5=(0)
          9'b010111100:  DATA = 16'b0000000000001000;    // h189_5=(0.00024414)
          9'b010111101:  DATA = 16'b0000000000001111;    // h190_5=(0.00045776)
          9'b010111110:  DATA = 16'b0000000000010111;    // h191_5=(0.0007019)
          9'b010111111:  DATA = 16'b0000000000011110;    // h192_5=(0.00091553)
          9'b011000000:  DATA = 16'b0000000000100110;    // h193_5=(0.0011597)
          9'b011000001:  DATA = 16'b0000000000101101;    // h194_5=(0.0013733)
          9'b011000010:  DATA = 16'b0000000000110100;    // h195_5=(0.0015869)
          9'b011000011:  DATA = 16'b0000000000111011;    // h196_5=(0.0018005)
          9'b011000100:  DATA = 16'b0000000001000010;    // h197_5=(0.0020142)
          9'b011000101:  DATA = 16'b0000000001001001;    // h198_5=(0.0022278)
          9'b011000110:  DATA = 16'b0000000001001111;    // h199_5=(0.0024109)
          9'b011000111:  DATA = 16'b0000000001010110;    // h200_5=(0.0026245)
          9'b011001000:  DATA = 16'b0000000001011101;    // h201_5=(0.0028381)
          9'b011001001:  DATA = 16'b0000000001100011;    // h202_5=(0.0030212)
          9'b011001010:  DATA = 16'b0000000001101001;    // h203_5=(0.0032043)
          9'b011001011:  DATA = 16'b0000000001101111;    // h204_5=(0.0033875)
          9'b011001100:  DATA = 16'b0000000001110101;    // h205_5=(0.0035706)
          9'b011001101:  DATA = 16'b0000000001111011;    // h206_5=(0.0037537)
          9'b011001110:  DATA = 16'b0000000010000001;    // h207_5=(0.0039368)
          9'b011001111:  DATA = 16'b0000000010000111;    // h208_5=(0.0041199)
          9'b011010000:  DATA = 16'b0000000010001100;    // h209_5=(0.0042725)
          9'b011010001:  DATA = 16'b0000000010010010;    // h210_5=(0.0044556)
          9'b011010010:  DATA = 16'b0000000010010111;    // h211_5=(0.0046082)
          9'b011010011:  DATA = 16'b0000000010011101;    // h212_5=(0.0047913)
          9'b011010100:  DATA = 16'b0000000010100010;    // h213_5=(0.0049438)
          9'b011010101:  DATA = 16'b0000000010100111;    // h214_5=(0.0050964)
          9'b011010110:  DATA = 16'b0000000010101100;    // h215_5=(0.005249)
          9'b011010111:  DATA = 16'b0000000010110001;    // h216_5=(0.0054016)
          9'b011011000:  DATA = 16'b0000000010110110;    // h217_5=(0.0055542)
          9'b011011001:  DATA = 16'b0000000010111010;    // h218_5=(0.0056763)
          9'b011011010:  DATA = 16'b0000000010111111;    // h219_5=(0.0058289)
          9'b011011011:  DATA = 16'b0000000011000100;    // h220_5=(0.0059814)
          9'b011011100:  DATA = 16'b0000000011001000;    // h221_5=(0.0061035)
          9'b011011101:  DATA = 16'b0000000011001100;    // h222_5=(0.0062256)
          9'b011011110:  DATA = 16'b0000000011010001;    // h223_5=(0.0063782)
          9'b011011111:  DATA = 16'b0000000011010101;    // h224_5=(0.0065002)
          9'b011100000:  DATA = 16'b0000000011011001;    // h225_5=(0.0066223)
          9'b011100001:  DATA = 16'b0000000011011101;    // h226_5=(0.0067444)
          9'b011100010:  DATA = 16'b0000000011100000;    // h227_5=(0.0068359)
          9'b011100011:  DATA = 16'b0000000011100100;    // h228_5=(0.006958)
          9'b011100100:  DATA = 16'b0000000011101000;    // h229_5=(0.0070801)
          9'b011100101:  DATA = 16'b0000000011101011;    // h230_5=(0.0071716)
          9'b011100110:  DATA = 16'b0000000011101111;    // h231_5=(0.0072937)
          9'b011100111:  DATA = 16'b0000000011110010;    // h232_5=(0.0073853)
          9'b011101000:  DATA = 16'b0000000011110110;    // h233_5=(0.0075073)
          9'b011101001:  DATA = 16'b0000000011111001;    // h234_5=(0.0075989)
          9'b011101010:  DATA = 16'b0000000011111100;    // h235_5=(0.0076904)
          9'b011101011:  DATA = 16'b0000000011111111;    // h236_5=(0.007782)
          9'b011101100:  DATA = 16'b0000000100000010;    // h237_5=(0.0078735)
          9'b011101101:  DATA = 16'b0000000100000101;    // h238_5=(0.0079651)
          9'b011101110:  DATA = 16'b0000000100001000;    // h239_5=(0.0080566)
          9'b011101111:  DATA = 16'b0000000100001010;    // h240_5=(0.0081177)
          9'b011110000:  DATA = 16'b0000000100001101;    // h241_5=(0.0082092)
          9'b011110001:  DATA = 16'b0000000100001111;    // h242_5=(0.0082703)
          9'b011110010:  DATA = 16'b0000000100010010;    // h243_5=(0.0083618)
          9'b011110011:  DATA = 16'b0000000100010100;    // h244_5=(0.0084229)
          9'b011110100:  DATA = 16'b0000000100010110;    // h245_5=(0.0084839)
          9'b011110101:  DATA = 16'b0000000100011001;    // h246_5=(0.0085754)
          9'b011110110:  DATA = 16'b0000000100011011;    // h247_5=(0.0086365)
          9'b011110111:  DATA = 16'b0000000100011101;    // h248_5=(0.0086975)
          9'b011111000:  DATA = 16'b0000000100011111;    // h249_5=(0.0087585)
          9'b011111001:  DATA = 16'b0000000100100000;    // h250_5=(0.0087891)
          9'b011111010:  DATA = 16'b0000000100100010;    // h251_5=(0.0088501)
          9'b011111011:  DATA = 16'b0000000100100100;    // h252_5=(0.0089111)
          9'b011111100:  DATA = 16'b0000000100100110;    // h253_5=(0.0089722)
          9'b011111101:  DATA = 16'b0000000100100111;    // h254_5=(0.0090027)
          9'b011111110:  DATA = 16'b0000000100101001;    // h255_5=(0.0090637)
          9'b011111111:  DATA = 16'b0000000100101010;    // h256_5=(0.0090942)
          9'b100000000:  DATA = 16'b0000000100101011;    // h257_5=(0.0091248)
          9'b100000001:  DATA = 16'b0000000100101101;    // h258_5=(0.0091858)
          9'b100000010:  DATA = 16'b0000000100101110;    // h259_5=(0.0092163)
          9'b100000011:  DATA = 16'b0000000100101111;    // h260_5=(0.0092468)
          9'b100000100:  DATA = 16'b0000000100110000;    // h261_5=(0.0092773)
          9'b100000101:  DATA = 16'b0000000100110001;    // h262_5=(0.0093079)
          9'b100000110:  DATA = 16'b0000000100110010;    // h263_5=(0.0093384)
          9'b100000111:  DATA = 16'b0000000100110011;    // h264_5=(0.0093689)
          9'b100001000:  DATA = 16'b0000000100110100;    // h265_5=(0.0093994)
          9'b100001001:  DATA = 16'b0000000100110100;    // h266_5=(0.0093994)
          9'b100001010:  DATA = 16'b0000000100110101;    // h267_5=(0.0094299)
          9'b100001011:  DATA = 16'b0000000100110110;    // h268_5=(0.0094604)
          9'b100001100:  DATA = 16'b0000000100110110;    // h269_5=(0.0094604)
          9'b100001101:  DATA = 16'b0000000100110111;    // h270_5=(0.009491)
          9'b100001110:  DATA = 16'b0000000100110111;    // h271_5=(0.009491)
          9'b100001111:  DATA = 16'b0000000100110111;    // h272_5=(0.009491)
          9'b100010000:  DATA = 16'b0000000100111000;    // h273_5=(0.0095215)
          9'b100010001:  DATA = 16'b0000000100111000;    // h274_5=(0.0095215)
          9'b100010010:  DATA = 16'b0000000100111000;    // h275_5=(0.0095215)
          9'b100010011:  DATA = 16'b0000000100111000;    // h276_5=(0.0095215)
          9'b100010100:  DATA = 16'b0000000100111000;    // h277_5=(0.0095215)
          9'b100010101:  DATA = 16'b0000000100111000;    // h278_5=(0.0095215)
          9'b100010110:  DATA = 16'b0000000100111000;    // h279_5=(0.0095215)
          9'b100010111:  DATA = 16'b0000000100111000;    // h280_5=(0.0095215)
          9'b100011000:  DATA = 16'b0000000100111000;    // h281_5=(0.0095215)
          9'b100011001:  DATA = 16'b0000000100110111;    // h282_5=(0.009491)
          9'b100011010:  DATA = 16'b0000000100110111;    // h283_5=(0.009491)
          9'b100011011:  DATA = 16'b0000000100110111;    // h284_5=(0.009491)
          9'b100011100:  DATA = 16'b0000000100110110;    // h285_5=(0.0094604)
          9'b100011101:  DATA = 16'b0000000100110110;    // h286_5=(0.0094604)
          9'b100011110:  DATA = 16'b0000000100110101;    // h287_5=(0.0094299)
          9'b100011111:  DATA = 16'b0000000100110101;    // h288_5=(0.0094299)
          9'b100100000:  DATA = 16'b0000000100110100;    // h289_5=(0.0093994)
          9'b100100001:  DATA = 16'b0000000100110100;    // h290_5=(0.0093994)
          9'b100100010:  DATA = 16'b0000000100110011;    // h291_5=(0.0093689)
          9'b100100011:  DATA = 16'b0000000100110010;    // h292_5=(0.0093384)
          9'b100100100:  DATA = 16'b0000000100110001;    // h293_5=(0.0093079)
          9'b100100101:  DATA = 16'b0000000100110001;    // h294_5=(0.0093079)
          9'b100100110:  DATA = 16'b0000000100110000;    // h295_5=(0.0092773)
          9'b100100111:  DATA = 16'b0000000100101111;    // h296_5=(0.0092468)
          9'b100101000:  DATA = 16'b0000000100101110;    // h297_5=(0.0092163)
          9'b100101001:  DATA = 16'b0000000100101101;    // h298_5=(0.0091858)
          9'b100101010:  DATA = 16'b0000000100101100;    // h299_5=(0.0091553)
          9'b100101011:  DATA = 16'b0000000100101011;    // h300_5=(0.0091248)
          9'b100101100:  DATA = 16'b0000000100101010;    // h301_5=(0.0090942)
          9'b100101101:  DATA = 16'b0000000100101000;    // h302_5=(0.0090332)
          9'b100101110:  DATA = 16'b0000000100100111;    // h303_5=(0.0090027)
          9'b100101111:  DATA = 16'b0000000100100110;    // h304_5=(0.0089722)
          9'b100110000:  DATA = 16'b0000000100100101;    // h305_5=(0.0089417)
          9'b100110001:  DATA = 16'b0000000100100011;    // h306_5=(0.0088806)
          9'b100110010:  DATA = 16'b0000000100100010;    // h307_5=(0.0088501)
          9'b100110011:  DATA = 16'b0000000100100001;    // h308_5=(0.0088196)
          9'b100110100:  DATA = 16'b0000000100011111;    // h309_5=(0.0087585)
          9'b100110101:  DATA = 16'b0000000100011110;    // h310_5=(0.008728)
          9'b100110110:  DATA = 16'b0000000100011100;    // h311_5=(0.008667)
          9'b100110111:  DATA = 16'b0000000100011011;    // h312_5=(0.0086365)
          9'b100111000:  DATA = 16'b0000000100011001;    // h313_5=(0.0085754)
          9'b100111001:  DATA = 16'b0000000100011000;    // h314_5=(0.0085449)
          9'b100111010:  DATA = 16'b0000000100010110;    // h315_5=(0.0084839)
          9'b100111011:  DATA = 16'b0000000100010101;    // h316_5=(0.0084534)
          9'b100111100:  DATA = 16'b0000000100010011;    // h317_5=(0.0083923)
          9'b100111101:  DATA = 16'b0000000100010001;    // h318_5=(0.0083313)
          9'b100111110:  DATA = 16'b0000000100010000;    // h319_5=(0.0083008)
          9'b100111111:  DATA = 16'b0000000100001110;    // h320_5=(0.0082397)
          9'b101000000:  DATA = 16'b0000000100001100;    // h321_5=(0.0081787)
          9'b101000001:  DATA = 16'b0000000100001010;    // h322_5=(0.0081177)
          9'b101000010:  DATA = 16'b0000000100001001;    // h323_5=(0.0080872)
          9'b101000011:  DATA = 16'b0000000100000111;    // h324_5=(0.0080261)
          9'b101000100:  DATA = 16'b0000000100000101;    // h325_5=(0.0079651)
          9'b101000101:  DATA = 16'b0000000100000011;    // h326_5=(0.0079041)
          9'b101000110:  DATA = 16'b0000000100000001;    // h327_5=(0.007843)
          9'b101000111:  DATA = 16'b0000000011111111;    // h328_5=(0.007782)
          9'b101001000:  DATA = 16'b0000000011111101;    // h329_5=(0.0077209)
          9'b101001001:  DATA = 16'b0000000011111011;    // h330_5=(0.0076599)
          9'b101001010:  DATA = 16'b0000000011111001;    // h331_5=(0.0075989)
          9'b101001011:  DATA = 16'b0000000011110111;    // h332_5=(0.0075378)
          9'b101001100:  DATA = 16'b0000000011110101;    // h333_5=(0.0074768)
          9'b101001101:  DATA = 16'b0000000011110011;    // h334_5=(0.0074158)
          9'b101001110:  DATA = 16'b0000000011110001;    // h335_5=(0.0073547)
          9'b101001111:  DATA = 16'b0000000011101111;    // h336_5=(0.0072937)
          9'b101010000:  DATA = 16'b0000000011101101;    // h337_5=(0.0072327)
          9'b101010001:  DATA = 16'b0000000011101011;    // h338_5=(0.0071716)
          9'b101010010:  DATA = 16'b0000000011101001;    // h339_5=(0.0071106)
          9'b101010011:  DATA = 16'b0000000011100111;    // h340_5=(0.0070496)
          9'b101010100:  DATA = 16'b0000000011100101;    // h341_5=(0.0069885)
          9'b101010101:  DATA = 16'b0000000011100011;    // h342_5=(0.0069275)
          9'b101010110:  DATA = 16'b0000000011100001;    // h343_5=(0.0068665)
          9'b101010111:  DATA = 16'b0000000011011110;    // h344_5=(0.0067749)
          9'b101011000:  DATA = 16'b0000000011011100;    // h345_5=(0.0067139)
          9'b101011001:  DATA = 16'b0000000011011010;    // h346_5=(0.0066528)
          9'b101011010:  DATA = 16'b0000000011011000;    // h347_5=(0.0065918)
          9'b101011011:  DATA = 16'b0000000011010110;    // h348_5=(0.0065308)
          9'b101011100:  DATA = 16'b0000000011010100;    // h349_5=(0.0064697)
          9'b101011101:  DATA = 16'b0000000011010001;    // h350_5=(0.0063782)
          9'b101011110:  DATA = 16'b0000000011001111;    // h351_5=(0.0063171)
          9'b101011111:  DATA = 16'b0000000011001101;    // h352_5=(0.0062561)
          9'b101100000:  DATA = 16'b0000000011001011;    // h353_5=(0.0061951)
          9'b101100001:  DATA = 16'b0000000011001001;    // h354_5=(0.006134)
          9'b101100010:  DATA = 16'b0000000011000110;    // h355_5=(0.0060425)
          9'b101100011:  DATA = 16'b0000000011000100;    // h356_5=(0.0059814)
          9'b101100100:  DATA = 16'b0000000011000010;    // h357_5=(0.0059204)
          9'b101100101:  DATA = 16'b0000000011000000;    // h358_5=(0.0058594)
          9'b101100110:  DATA = 16'b0000000010111101;    // h359_5=(0.0057678)
          9'b101100111:  DATA = 16'b0000000010111011;    // h360_5=(0.0057068)
          9'b101101000:  DATA = 16'b0000000010111001;    // h361_5=(0.0056458)
          9'b101101001:  DATA = 16'b0000000010110111;    // h362_5=(0.0055847)
          9'b101101010:  DATA = 16'b0000000010110100;    // h363_5=(0.0054932)
          9'b101101011:  DATA = 16'b0000000010110010;    // h364_5=(0.0054321)
          9'b101101100:  DATA = 16'b0000000010110000;    // h365_5=(0.0053711)
          9'b101101101:  DATA = 16'b0000000010101110;    // h366_5=(0.0053101)
          9'b101101110:  DATA = 16'b0000000010101011;    // h367_5=(0.0052185)
          9'b101101111:  DATA = 16'b0000000010101001;    // h368_5=(0.0051575)
          9'b101110000:  DATA = 16'b0000000010100111;    // h369_5=(0.0050964)
          9'b101110001:  DATA = 16'b0000000010100101;    // h370_5=(0.0050354)
          9'b101110010:  DATA = 16'b0000000010100011;    // h371_5=(0.0049744)
          9'b101110011:  DATA = 16'b0000000010100000;    // h372_5=(0.0048828)
          9'b101110100:  DATA = 16'b0000000010011110;    // h373_5=(0.0048218)
          9'b101110101:  DATA = 16'b0000000010011100;    // h374_5=(0.0047607)
          9'b101110110:  DATA = 16'b0000000010011010;    // h375_5=(0.0046997)
          default : DATA = 16'b0000000000000000;
        endcase
    end
endmodule

