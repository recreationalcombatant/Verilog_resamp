`timescale 1ns / 1ps
///////////////////////////////////////////
// ROM table - 2's complement coefficients
// fir_rom3.v: FIR polyphase branch (3)
// 
// Created: 03-Aug-2006 17:33:00
//  from Matlab script fpga_create_rom_verilog.m
//
// J. Shima
//////////////////////////////////////////
module fir_rom3(ADDR, DATA);
    input [8:0] ADDR;
    output signed [15:0] DATA;
    reg signed [15:0] DATA;

    always@(ADDR) begin
        case(ADDR)
          9'b000000000:  DATA = 16'b0100101011100110;    // h1_3=(0.58514)
          9'b000000001:  DATA = 16'b0100101101011111;    // h2_3=(0.58884)
          9'b000000010:  DATA = 16'b0100101111010111;    // h3_3=(0.5925)
          9'b000000011:  DATA = 16'b0100110001001111;    // h4_3=(0.59616)
          9'b000000100:  DATA = 16'b0100110011000111;    // h5_3=(0.59982)
          9'b000000101:  DATA = 16'b0100110100111111;    // h6_3=(0.60349)
          9'b000000110:  DATA = 16'b0100110110110110;    // h7_3=(0.60712)
          9'b000000111:  DATA = 16'b0100111000101101;    // h8_3=(0.61075)
          9'b000001000:  DATA = 16'b0100111010100101;    // h9_3=(0.61441)
          9'b000001001:  DATA = 16'b0100111100011100;    // h10_3=(0.61804)
          9'b000001010:  DATA = 16'b0100111110010010;    // h11_3=(0.62164)
          9'b000001011:  DATA = 16'b0101000000001001;    // h12_3=(0.62527)
          9'b000001100:  DATA = 16'b0101000001111111;    // h13_3=(0.62888)
          9'b000001101:  DATA = 16'b0101000011110101;    // h14_3=(0.63248)
          9'b000001110:  DATA = 16'b0101000101101011;    // h15_3=(0.63608)
          9'b000001111:  DATA = 16'b0101000111100001;    // h16_3=(0.63968)
          9'b000010000:  DATA = 16'b0101001001010110;    // h17_3=(0.64325)
          9'b000010001:  DATA = 16'b0101001011001100;    // h18_3=(0.64685)
          9'b000010010:  DATA = 16'b0101001101000001;    // h19_3=(0.65042)
          9'b000010011:  DATA = 16'b0101001110110101;    // h20_3=(0.65396)
          9'b000010100:  DATA = 16'b0101010000101010;    // h21_3=(0.65753)
          9'b000010101:  DATA = 16'b0101010010011110;    // h22_3=(0.66107)
          9'b000010110:  DATA = 16'b0101010100010010;    // h23_3=(0.66461)
          9'b000010111:  DATA = 16'b0101010110000101;    // h24_3=(0.66812)
          9'b000011000:  DATA = 16'b0101010111111000;    // h25_3=(0.67163)
          9'b000011001:  DATA = 16'b0101011001101011;    // h26_3=(0.67514)
          9'b000011010:  DATA = 16'b0101011011011110;    // h27_3=(0.67865)
          9'b000011011:  DATA = 16'b0101011101010001;    // h28_3=(0.68216)
          9'b000011100:  DATA = 16'b0101011111000011;    // h29_3=(0.68564)
          9'b000011101:  DATA = 16'b0101100000110100;    // h30_3=(0.68909)
          9'b000011110:  DATA = 16'b0101100010100110;    // h31_3=(0.69257)
          9'b000011111:  DATA = 16'b0101100100010111;    // h32_3=(0.69601)
          9'b000100000:  DATA = 16'b0101100110000111;    // h33_3=(0.69943)
          9'b000100001:  DATA = 16'b0101100111111000;    // h34_3=(0.70288)
          9'b000100010:  DATA = 16'b0101101001101000;    // h35_3=(0.7063)
          9'b000100011:  DATA = 16'b0101101011011000;    // h36_3=(0.70972)
          9'b000100100:  DATA = 16'b0101101101000111;    // h37_3=(0.7131)
          9'b000100101:  DATA = 16'b0101101110110110;    // h38_3=(0.71649)
          9'b000100110:  DATA = 16'b0101110000100100;    // h39_3=(0.71985)
          9'b000100111:  DATA = 16'b0101110010010010;    // h40_3=(0.72321)
          9'b000101000:  DATA = 16'b0101110100000000;    // h41_3=(0.72656)
          9'b000101001:  DATA = 16'b0101110101101110;    // h42_3=(0.72992)
          9'b000101010:  DATA = 16'b0101110111011011;    // h43_3=(0.73325)
          9'b000101011:  DATA = 16'b0101111001000111;    // h44_3=(0.73654)
          9'b000101100:  DATA = 16'b0101111010110011;    // h45_3=(0.73984)
          9'b000101101:  DATA = 16'b0101111100011111;    // h46_3=(0.74313)
          9'b000101110:  DATA = 16'b0101111110001010;    // h47_3=(0.7464)
          9'b000101111:  DATA = 16'b0101111111110101;    // h48_3=(0.74966)
          9'b000110000:  DATA = 16'b0110000001011111;    // h49_3=(0.7529)
          9'b000110001:  DATA = 16'b0110000011001001;    // h50_3=(0.75613)
          9'b000110010:  DATA = 16'b0110000100110011;    // h51_3=(0.75937)
          9'b000110011:  DATA = 16'b0110000110011100;    // h52_3=(0.76257)
          9'b000110100:  DATA = 16'b0110001000000101;    // h53_3=(0.76578)
          9'b000110101:  DATA = 16'b0110001001101101;    // h54_3=(0.76895)
          9'b000110110:  DATA = 16'b0110001011010100;    // h55_3=(0.77209)
          9'b000110111:  DATA = 16'b0110001100111011;    // h56_3=(0.77524)
          9'b000111000:  DATA = 16'b0110001110100010;    // h57_3=(0.77838)
          9'b000111001:  DATA = 16'b0110010000001000;    // h58_3=(0.78149)
          9'b000111010:  DATA = 16'b0110010001101110;    // h59_3=(0.78461)
          9'b000111011:  DATA = 16'b0110010011010011;    // h60_3=(0.78769)
          9'b000111100:  DATA = 16'b0110010100111000;    // h61_3=(0.79077)
          9'b000111101:  DATA = 16'b0110010110011100;    // h62_3=(0.79382)
          9'b000111110:  DATA = 16'b0110010111111111;    // h63_3=(0.79684)
          9'b000111111:  DATA = 16'b0110011001100010;    // h64_3=(0.79987)
          9'b001000000:  DATA = 16'b0110011011000101;    // h65_3=(0.80289)
          9'b001000001:  DATA = 16'b0110011100100111;    // h66_3=(0.80588)
          9'b001000010:  DATA = 16'b0110011110001000;    // h67_3=(0.80884)
          9'b001000011:  DATA = 16'b0110011111101001;    // h68_3=(0.8118)
          9'b001000100:  DATA = 16'b0110100001001010;    // h69_3=(0.81476)
          9'b001000101:  DATA = 16'b0110100010101001;    // h70_3=(0.81766)
          9'b001000110:  DATA = 16'b0110100100001001;    // h71_3=(0.82059)
          9'b001000111:  DATA = 16'b0110100101100111;    // h72_3=(0.82346)
          9'b001001000:  DATA = 16'b0110100111000101;    // h73_3=(0.82632)
          9'b001001001:  DATA = 16'b0110101000100011;    // h74_3=(0.82919)
          9'b001001010:  DATA = 16'b0110101010000000;    // h75_3=(0.83203)
          9'b001001011:  DATA = 16'b0110101011011100;    // h76_3=(0.83484)
          9'b001001100:  DATA = 16'b0110101100110111;    // h77_3=(0.83762)
          9'b001001101:  DATA = 16'b0110101110010011;    // h78_3=(0.84042)
          9'b001001110:  DATA = 16'b0110101111101101;    // h79_3=(0.84317)
          9'b001001111:  DATA = 16'b0110110001000111;    // h80_3=(0.84592)
          9'b001010000:  DATA = 16'b0110110010100000;    // h81_3=(0.84863)
          9'b001010001:  DATA = 16'b0110110011111001;    // h82_3=(0.85135)
          9'b001010010:  DATA = 16'b0110110101010000;    // h83_3=(0.854)
          9'b001010011:  DATA = 16'b0110110110101000;    // h84_3=(0.85669)
          9'b001010100:  DATA = 16'b0110110111111110;    // h85_3=(0.85931)
          9'b001010101:  DATA = 16'b0110111001010100;    // h86_3=(0.86194)
          9'b001010110:  DATA = 16'b0110111010101010;    // h87_3=(0.86456)
          9'b001010111:  DATA = 16'b0110111011111110;    // h88_3=(0.86713)
          9'b001011000:  DATA = 16'b0110111101010010;    // h89_3=(0.86969)
          9'b001011001:  DATA = 16'b0110111110100110;    // h90_3=(0.87225)
          9'b001011010:  DATA = 16'b0110111111111000;    // h91_3=(0.87476)
          9'b001011011:  DATA = 16'b0111000001001010;    // h92_3=(0.87726)
          9'b001011100:  DATA = 16'b0111000010011100;    // h93_3=(0.87976)
          9'b001011101:  DATA = 16'b0111000011101100;    // h94_3=(0.8822)
          9'b001011110:  DATA = 16'b0111000100111100;    // h95_3=(0.88464)
          9'b001011111:  DATA = 16'b0111000110001011;    // h96_3=(0.88705)
          9'b001100000:  DATA = 16'b0111000111011010;    // h97_3=(0.88947)
          9'b001100001:  DATA = 16'b0111001000101000;    // h98_3=(0.89185)
          9'b001100010:  DATA = 16'b0111001001110101;    // h99_3=(0.8942)
          9'b001100011:  DATA = 16'b0111001011000001;    // h100_3=(0.89651)
          9'b001100100:  DATA = 16'b0111001100001101;    // h101_3=(0.89883)
          9'b001100101:  DATA = 16'b0111001101011000;    // h102_3=(0.90112)
          9'b001100110:  DATA = 16'b0111001110100010;    // h103_3=(0.90338)
          9'b001100111:  DATA = 16'b0111001111101011;    // h104_3=(0.90561)
          9'b001101000:  DATA = 16'b0111010000110100;    // h105_3=(0.90784)
          9'b001101001:  DATA = 16'b0111010001111100;    // h106_3=(0.91003)
          9'b001101010:  DATA = 16'b0111010011000011;    // h107_3=(0.9122)
          9'b001101011:  DATA = 16'b0111010100001001;    // h108_3=(0.91434)
          9'b001101100:  DATA = 16'b0111010101001111;    // h109_3=(0.91647)
          9'b001101101:  DATA = 16'b0111010110010100;    // h110_3=(0.91858)
          9'b001101110:  DATA = 16'b0111010111011000;    // h111_3=(0.92065)
          9'b001101111:  DATA = 16'b0111011000011100;    // h112_3=(0.92273)
          9'b001110000:  DATA = 16'b0111011001011110;    // h113_3=(0.92474)
          9'b001110001:  DATA = 16'b0111011010100000;    // h114_3=(0.92676)
          9'b001110010:  DATA = 16'b0111011011100001;    // h115_3=(0.92874)
          9'b001110011:  DATA = 16'b0111011100100001;    // h116_3=(0.93069)
          9'b001110100:  DATA = 16'b0111011101100001;    // h117_3=(0.93265)
          9'b001110101:  DATA = 16'b0111011110011111;    // h118_3=(0.93454)
          9'b001110110:  DATA = 16'b0111011111011101;    // h119_3=(0.93643)
          9'b001110111:  DATA = 16'b0111100000011010;    // h120_3=(0.93829)
          9'b001111000:  DATA = 16'b0111100001010111;    // h121_3=(0.94016)
          9'b001111001:  DATA = 16'b0111100010010010;    // h122_3=(0.94196)
          9'b001111010:  DATA = 16'b0111100011001101;    // h123_3=(0.94376)
          9'b001111011:  DATA = 16'b0111100100000111;    // h124_3=(0.94553)
          9'b001111100:  DATA = 16'b0111100101000000;    // h125_3=(0.94727)
          9'b001111101:  DATA = 16'b0111100101111000;    // h126_3=(0.94897)
          9'b001111110:  DATA = 16'b0111100110101111;    // h127_3=(0.95065)
          9'b001111111:  DATA = 16'b0111100111100110;    // h128_3=(0.95233)
          9'b010000000:  DATA = 16'b0111101000011011;    // h129_3=(0.95395)
          9'b010000001:  DATA = 16'b0111101001010000;    // h130_3=(0.95557)
          9'b010000010:  DATA = 16'b0111101010000100;    // h131_3=(0.95715)
          9'b010000011:  DATA = 16'b0111101010110111;    // h132_3=(0.95871)
          9'b010000100:  DATA = 16'b0111101011101010;    // h133_3=(0.96027)
          9'b010000101:  DATA = 16'b0111101100011011;    // h134_3=(0.96176)
          9'b010000110:  DATA = 16'b0111101101001100;    // h135_3=(0.96326)
          9'b010000111:  DATA = 16'b0111101101111011;    // h136_3=(0.96469)
          9'b010001000:  DATA = 16'b0111101110101010;    // h137_3=(0.96613)
          9'b010001001:  DATA = 16'b0111101111011000;    // h138_3=(0.96753)
          9'b010001010:  DATA = 16'b0111110000000110;    // h139_3=(0.96893)
          9'b010001011:  DATA = 16'b0111110000110010;    // h140_3=(0.97028)
          9'b010001100:  DATA = 16'b0111110001011101;    // h141_3=(0.97159)
          9'b010001101:  DATA = 16'b0111110010001000;    // h142_3=(0.9729)
          9'b010001110:  DATA = 16'b0111110010110010;    // h143_3=(0.97418)
          9'b010001111:  DATA = 16'b0111110011011010;    // h144_3=(0.9754)
          9'b010010000:  DATA = 16'b0111110100000010;    // h145_3=(0.97662)
          9'b010010001:  DATA = 16'b0111110100101001;    // h146_3=(0.97781)
          9'b010010010:  DATA = 16'b0111110101001111;    // h147_3=(0.97897)
          9'b010010011:  DATA = 16'b0111110101110101;    // h148_3=(0.98013)
          9'b010010100:  DATA = 16'b0111110110011001;    // h149_3=(0.98123)
          9'b010010101:  DATA = 16'b0111110110111101;    // h150_3=(0.98233)
          9'b010010110:  DATA = 16'b0111110111011111;    // h151_3=(0.98337)
          9'b010010111:  DATA = 16'b0111111000000001;    // h152_3=(0.98441)
          9'b010011000:  DATA = 16'b0111111000100010;    // h153_3=(0.98541)
          9'b010011001:  DATA = 16'b0111111001000010;    // h154_3=(0.98639)
          9'b010011010:  DATA = 16'b0111111001100001;    // h155_3=(0.98734)
          9'b010011011:  DATA = 16'b0111111001111111;    // h156_3=(0.98825)
          9'b010011100:  DATA = 16'b0111111010011100;    // h157_3=(0.98914)
          9'b010011101:  DATA = 16'b0111111010111000;    // h158_3=(0.98999)
          9'b010011110:  DATA = 16'b0111111011010011;    // h159_3=(0.99081)
          9'b010011111:  DATA = 16'b0111111011101110;    // h160_3=(0.99164)
          9'b010100000:  DATA = 16'b0111111100000111;    // h161_3=(0.9924)
          9'b010100001:  DATA = 16'b0111111100100000;    // h162_3=(0.99316)
          9'b010100010:  DATA = 16'b0111111100111000;    // h163_3=(0.9939)
          9'b010100011:  DATA = 16'b0111111101001111;    // h164_3=(0.9946)
          9'b010100100:  DATA = 16'b0111111101100100;    // h165_3=(0.99524)
          9'b010100101:  DATA = 16'b0111111101111001;    // h166_3=(0.99588)
          9'b010100110:  DATA = 16'b0111111110001101;    // h167_3=(0.99649)
          9'b010100111:  DATA = 16'b0111111110100001;    // h168_3=(0.9971)
          9'b010101000:  DATA = 16'b0111111110110011;    // h169_3=(0.99765)
          9'b010101001:  DATA = 16'b0111111111000100;    // h170_3=(0.99817)
          9'b010101010:  DATA = 16'b0111111111010100;    // h171_3=(0.99866)
          9'b010101011:  DATA = 16'b0111111111100100;    // h172_3=(0.99915)
          9'b010101100:  DATA = 16'b0111111111110010;    // h173_3=(0.99957)
          9'b010101101:  DATA = 16'b0111111111111111;    // h174_3=(0.99997)
          9'b010101110:  DATA = 16'b0111111111111111;    // h175_3=(0.99997)
          9'b010101111:  DATA = 16'b0111111111111111;    // h176_3=(0.99997)
          9'b010110000:  DATA = 16'b0111111111111111;    // h177_3=(0.99997)
          9'b010110001:  DATA = 16'b0111111111111111;    // h178_3=(0.99997)
          9'b010110010:  DATA = 16'b0111111111111111;    // h179_3=(0.99997)
          9'b010110011:  DATA = 16'b0111111111111111;    // h180_3=(0.99997)
          9'b010110100:  DATA = 16'b0111111111111111;    // h181_3=(0.99997)
          9'b010110101:  DATA = 16'b0111111111111111;    // h182_3=(0.99997)
          9'b010110110:  DATA = 16'b0111111111111111;    // h183_3=(0.99997)
          9'b010110111:  DATA = 16'b0111111111111111;    // h184_3=(0.99997)
          9'b010111000:  DATA = 16'b0111111111111111;    // h185_3=(0.99997)
          9'b010111001:  DATA = 16'b0111111111111111;    // h186_3=(0.99997)
          9'b010111010:  DATA = 16'b0111111111111111;    // h187_3=(0.99997)
          9'b010111011:  DATA = 16'b0111111111111111;    // h188_3=(0.99997)
          9'b010111100:  DATA = 16'b0111111111111111;    // h189_3=(0.99997)
          9'b010111101:  DATA = 16'b0111111111111111;    // h190_3=(0.99997)
          9'b010111110:  DATA = 16'b0111111111111111;    // h191_3=(0.99997)
          9'b010111111:  DATA = 16'b0111111111111111;    // h192_3=(0.99997)
          9'b011000000:  DATA = 16'b0111111111111111;    // h193_3=(0.99997)
          9'b011000001:  DATA = 16'b0111111111111111;    // h194_3=(0.99997)
          9'b011000010:  DATA = 16'b0111111111111111;    // h195_3=(0.99997)
          9'b011000011:  DATA = 16'b0111111111111111;    // h196_3=(0.99997)
          9'b011000100:  DATA = 16'b0111111111111111;    // h197_3=(0.99997)
          9'b011000101:  DATA = 16'b0111111111111111;    // h198_3=(0.99997)
          9'b011000110:  DATA = 16'b0111111111111111;    // h199_3=(0.99997)
          9'b011000111:  DATA = 16'b0111111111111111;    // h200_3=(0.99997)
          9'b011001000:  DATA = 16'b0111111111111111;    // h201_3=(0.99997)
          9'b011001001:  DATA = 16'b0111111111111111;    // h202_3=(0.99997)
          9'b011001010:  DATA = 16'b0111111111110010;    // h203_3=(0.99957)
          9'b011001011:  DATA = 16'b0111111111100100;    // h204_3=(0.99915)
          9'b011001100:  DATA = 16'b0111111111010100;    // h205_3=(0.99866)
          9'b011001101:  DATA = 16'b0111111111000100;    // h206_3=(0.99817)
          9'b011001110:  DATA = 16'b0111111110110011;    // h207_3=(0.99765)
          9'b011001111:  DATA = 16'b0111111110100001;    // h208_3=(0.9971)
          9'b011010000:  DATA = 16'b0111111110001101;    // h209_3=(0.99649)
          9'b011010001:  DATA = 16'b0111111101111001;    // h210_3=(0.99588)
          9'b011010010:  DATA = 16'b0111111101100100;    // h211_3=(0.99524)
          9'b011010011:  DATA = 16'b0111111101001111;    // h212_3=(0.9946)
          9'b011010100:  DATA = 16'b0111111100111000;    // h213_3=(0.9939)
          9'b011010101:  DATA = 16'b0111111100100000;    // h214_3=(0.99316)
          9'b011010110:  DATA = 16'b0111111100000111;    // h215_3=(0.9924)
          9'b011010111:  DATA = 16'b0111111011101110;    // h216_3=(0.99164)
          9'b011011000:  DATA = 16'b0111111011010011;    // h217_3=(0.99081)
          9'b011011001:  DATA = 16'b0111111010111000;    // h218_3=(0.98999)
          9'b011011010:  DATA = 16'b0111111010011100;    // h219_3=(0.98914)
          9'b011011011:  DATA = 16'b0111111001111111;    // h220_3=(0.98825)
          9'b011011100:  DATA = 16'b0111111001100001;    // h221_3=(0.98734)
          9'b011011101:  DATA = 16'b0111111001000010;    // h222_3=(0.98639)
          9'b011011110:  DATA = 16'b0111111000100010;    // h223_3=(0.98541)
          9'b011011111:  DATA = 16'b0111111000000001;    // h224_3=(0.98441)
          9'b011100000:  DATA = 16'b0111110111011111;    // h225_3=(0.98337)
          9'b011100001:  DATA = 16'b0111110110111101;    // h226_3=(0.98233)
          9'b011100010:  DATA = 16'b0111110110011001;    // h227_3=(0.98123)
          9'b011100011:  DATA = 16'b0111110101110101;    // h228_3=(0.98013)
          9'b011100100:  DATA = 16'b0111110101001111;    // h229_3=(0.97897)
          9'b011100101:  DATA = 16'b0111110100101001;    // h230_3=(0.97781)
          9'b011100110:  DATA = 16'b0111110100000010;    // h231_3=(0.97662)
          9'b011100111:  DATA = 16'b0111110011011010;    // h232_3=(0.9754)
          9'b011101000:  DATA = 16'b0111110010110010;    // h233_3=(0.97418)
          9'b011101001:  DATA = 16'b0111110010001000;    // h234_3=(0.9729)
          9'b011101010:  DATA = 16'b0111110001011101;    // h235_3=(0.97159)
          9'b011101011:  DATA = 16'b0111110000110010;    // h236_3=(0.97028)
          9'b011101100:  DATA = 16'b0111110000000110;    // h237_3=(0.96893)
          9'b011101101:  DATA = 16'b0111101111011000;    // h238_3=(0.96753)
          9'b011101110:  DATA = 16'b0111101110101010;    // h239_3=(0.96613)
          9'b011101111:  DATA = 16'b0111101101111011;    // h240_3=(0.96469)
          9'b011110000:  DATA = 16'b0111101101001100;    // h241_3=(0.96326)
          9'b011110001:  DATA = 16'b0111101100011011;    // h242_3=(0.96176)
          9'b011110010:  DATA = 16'b0111101011101010;    // h243_3=(0.96027)
          9'b011110011:  DATA = 16'b0111101010110111;    // h244_3=(0.95871)
          9'b011110100:  DATA = 16'b0111101010000100;    // h245_3=(0.95715)
          9'b011110101:  DATA = 16'b0111101001010000;    // h246_3=(0.95557)
          9'b011110110:  DATA = 16'b0111101000011011;    // h247_3=(0.95395)
          9'b011110111:  DATA = 16'b0111100111100110;    // h248_3=(0.95233)
          9'b011111000:  DATA = 16'b0111100110101111;    // h249_3=(0.95065)
          9'b011111001:  DATA = 16'b0111100101111000;    // h250_3=(0.94897)
          9'b011111010:  DATA = 16'b0111100101000000;    // h251_3=(0.94727)
          9'b011111011:  DATA = 16'b0111100100000111;    // h252_3=(0.94553)
          9'b011111100:  DATA = 16'b0111100011001101;    // h253_3=(0.94376)
          9'b011111101:  DATA = 16'b0111100010010010;    // h254_3=(0.94196)
          9'b011111110:  DATA = 16'b0111100001010111;    // h255_3=(0.94016)
          9'b011111111:  DATA = 16'b0111100000011010;    // h256_3=(0.93829)
          9'b100000000:  DATA = 16'b0111011111011101;    // h257_3=(0.93643)
          9'b100000001:  DATA = 16'b0111011110011111;    // h258_3=(0.93454)
          9'b100000010:  DATA = 16'b0111011101100001;    // h259_3=(0.93265)
          9'b100000011:  DATA = 16'b0111011100100001;    // h260_3=(0.93069)
          9'b100000100:  DATA = 16'b0111011011100001;    // h261_3=(0.92874)
          9'b100000101:  DATA = 16'b0111011010100000;    // h262_3=(0.92676)
          9'b100000110:  DATA = 16'b0111011001011110;    // h263_3=(0.92474)
          9'b100000111:  DATA = 16'b0111011000011100;    // h264_3=(0.92273)
          9'b100001000:  DATA = 16'b0111010111011000;    // h265_3=(0.92065)
          9'b100001001:  DATA = 16'b0111010110010100;    // h266_3=(0.91858)
          9'b100001010:  DATA = 16'b0111010101001111;    // h267_3=(0.91647)
          9'b100001011:  DATA = 16'b0111010100001001;    // h268_3=(0.91434)
          9'b100001100:  DATA = 16'b0111010011000011;    // h269_3=(0.9122)
          9'b100001101:  DATA = 16'b0111010001111100;    // h270_3=(0.91003)
          9'b100001110:  DATA = 16'b0111010000110100;    // h271_3=(0.90784)
          9'b100001111:  DATA = 16'b0111001111101011;    // h272_3=(0.90561)
          9'b100010000:  DATA = 16'b0111001110100010;    // h273_3=(0.90338)
          9'b100010001:  DATA = 16'b0111001101011000;    // h274_3=(0.90112)
          9'b100010010:  DATA = 16'b0111001100001101;    // h275_3=(0.89883)
          9'b100010011:  DATA = 16'b0111001011000001;    // h276_3=(0.89651)
          9'b100010100:  DATA = 16'b0111001001110101;    // h277_3=(0.8942)
          9'b100010101:  DATA = 16'b0111001000101000;    // h278_3=(0.89185)
          9'b100010110:  DATA = 16'b0111000111011010;    // h279_3=(0.88947)
          9'b100010111:  DATA = 16'b0111000110001011;    // h280_3=(0.88705)
          9'b100011000:  DATA = 16'b0111000100111100;    // h281_3=(0.88464)
          9'b100011001:  DATA = 16'b0111000011101100;    // h282_3=(0.8822)
          9'b100011010:  DATA = 16'b0111000010011100;    // h283_3=(0.87976)
          9'b100011011:  DATA = 16'b0111000001001010;    // h284_3=(0.87726)
          9'b100011100:  DATA = 16'b0110111111111000;    // h285_3=(0.87476)
          9'b100011101:  DATA = 16'b0110111110100110;    // h286_3=(0.87225)
          9'b100011110:  DATA = 16'b0110111101010010;    // h287_3=(0.86969)
          9'b100011111:  DATA = 16'b0110111011111110;    // h288_3=(0.86713)
          9'b100100000:  DATA = 16'b0110111010101010;    // h289_3=(0.86456)
          9'b100100001:  DATA = 16'b0110111001010100;    // h290_3=(0.86194)
          9'b100100010:  DATA = 16'b0110110111111110;    // h291_3=(0.85931)
          9'b100100011:  DATA = 16'b0110110110101000;    // h292_3=(0.85669)
          9'b100100100:  DATA = 16'b0110110101010000;    // h293_3=(0.854)
          9'b100100101:  DATA = 16'b0110110011111001;    // h294_3=(0.85135)
          9'b100100110:  DATA = 16'b0110110010100000;    // h295_3=(0.84863)
          9'b100100111:  DATA = 16'b0110110001000111;    // h296_3=(0.84592)
          9'b100101000:  DATA = 16'b0110101111101101;    // h297_3=(0.84317)
          9'b100101001:  DATA = 16'b0110101110010011;    // h298_3=(0.84042)
          9'b100101010:  DATA = 16'b0110101100110111;    // h299_3=(0.83762)
          9'b100101011:  DATA = 16'b0110101011011100;    // h300_3=(0.83484)
          9'b100101100:  DATA = 16'b0110101010000000;    // h301_3=(0.83203)
          9'b100101101:  DATA = 16'b0110101000100011;    // h302_3=(0.82919)
          9'b100101110:  DATA = 16'b0110100111000101;    // h303_3=(0.82632)
          9'b100101111:  DATA = 16'b0110100101100111;    // h304_3=(0.82346)
          9'b100110000:  DATA = 16'b0110100100001001;    // h305_3=(0.82059)
          9'b100110001:  DATA = 16'b0110100010101001;    // h306_3=(0.81766)
          9'b100110010:  DATA = 16'b0110100001001010;    // h307_3=(0.81476)
          9'b100110011:  DATA = 16'b0110011111101001;    // h308_3=(0.8118)
          9'b100110100:  DATA = 16'b0110011110001000;    // h309_3=(0.80884)
          9'b100110101:  DATA = 16'b0110011100100111;    // h310_3=(0.80588)
          9'b100110110:  DATA = 16'b0110011011000101;    // h311_3=(0.80289)
          9'b100110111:  DATA = 16'b0110011001100010;    // h312_3=(0.79987)
          9'b100111000:  DATA = 16'b0110010111111111;    // h313_3=(0.79684)
          9'b100111001:  DATA = 16'b0110010110011100;    // h314_3=(0.79382)
          9'b100111010:  DATA = 16'b0110010100111000;    // h315_3=(0.79077)
          9'b100111011:  DATA = 16'b0110010011010011;    // h316_3=(0.78769)
          9'b100111100:  DATA = 16'b0110010001101110;    // h317_3=(0.78461)
          9'b100111101:  DATA = 16'b0110010000001000;    // h318_3=(0.78149)
          9'b100111110:  DATA = 16'b0110001110100010;    // h319_3=(0.77838)
          9'b100111111:  DATA = 16'b0110001100111011;    // h320_3=(0.77524)
          9'b101000000:  DATA = 16'b0110001011010100;    // h321_3=(0.77209)
          9'b101000001:  DATA = 16'b0110001001101101;    // h322_3=(0.76895)
          9'b101000010:  DATA = 16'b0110001000000101;    // h323_3=(0.76578)
          9'b101000011:  DATA = 16'b0110000110011100;    // h324_3=(0.76257)
          9'b101000100:  DATA = 16'b0110000100110011;    // h325_3=(0.75937)
          9'b101000101:  DATA = 16'b0110000011001001;    // h326_3=(0.75613)
          9'b101000110:  DATA = 16'b0110000001011111;    // h327_3=(0.7529)
          9'b101000111:  DATA = 16'b0101111111110101;    // h328_3=(0.74966)
          9'b101001000:  DATA = 16'b0101111110001010;    // h329_3=(0.7464)
          9'b101001001:  DATA = 16'b0101111100011111;    // h330_3=(0.74313)
          9'b101001010:  DATA = 16'b0101111010110011;    // h331_3=(0.73984)
          9'b101001011:  DATA = 16'b0101111001000111;    // h332_3=(0.73654)
          9'b101001100:  DATA = 16'b0101110111011011;    // h333_3=(0.73325)
          9'b101001101:  DATA = 16'b0101110101101110;    // h334_3=(0.72992)
          9'b101001110:  DATA = 16'b0101110100000000;    // h335_3=(0.72656)
          9'b101001111:  DATA = 16'b0101110010010010;    // h336_3=(0.72321)
          9'b101010000:  DATA = 16'b0101110000100100;    // h337_3=(0.71985)
          9'b101010001:  DATA = 16'b0101101110110110;    // h338_3=(0.71649)
          9'b101010010:  DATA = 16'b0101101101000111;    // h339_3=(0.7131)
          9'b101010011:  DATA = 16'b0101101011011000;    // h340_3=(0.70972)
          9'b101010100:  DATA = 16'b0101101001101000;    // h341_3=(0.7063)
          9'b101010101:  DATA = 16'b0101100111111000;    // h342_3=(0.70288)
          9'b101010110:  DATA = 16'b0101100110000111;    // h343_3=(0.69943)
          9'b101010111:  DATA = 16'b0101100100010111;    // h344_3=(0.69601)
          9'b101011000:  DATA = 16'b0101100010100110;    // h345_3=(0.69257)
          9'b101011001:  DATA = 16'b0101100000110100;    // h346_3=(0.68909)
          9'b101011010:  DATA = 16'b0101011111000011;    // h347_3=(0.68564)
          9'b101011011:  DATA = 16'b0101011101010001;    // h348_3=(0.68216)
          9'b101011100:  DATA = 16'b0101011011011110;    // h349_3=(0.67865)
          9'b101011101:  DATA = 16'b0101011001101011;    // h350_3=(0.67514)
          9'b101011110:  DATA = 16'b0101010111111000;    // h351_3=(0.67163)
          9'b101011111:  DATA = 16'b0101010110000101;    // h352_3=(0.66812)
          9'b101100000:  DATA = 16'b0101010100010010;    // h353_3=(0.66461)
          9'b101100001:  DATA = 16'b0101010010011110;    // h354_3=(0.66107)
          9'b101100010:  DATA = 16'b0101010000101010;    // h355_3=(0.65753)
          9'b101100011:  DATA = 16'b0101001110110101;    // h356_3=(0.65396)
          9'b101100100:  DATA = 16'b0101001101000001;    // h357_3=(0.65042)
          9'b101100101:  DATA = 16'b0101001011001100;    // h358_3=(0.64685)
          9'b101100110:  DATA = 16'b0101001001010110;    // h359_3=(0.64325)
          9'b101100111:  DATA = 16'b0101000111100001;    // h360_3=(0.63968)
          9'b101101000:  DATA = 16'b0101000101101011;    // h361_3=(0.63608)
          9'b101101001:  DATA = 16'b0101000011110101;    // h362_3=(0.63248)
          9'b101101010:  DATA = 16'b0101000001111111;    // h363_3=(0.62888)
          9'b101101011:  DATA = 16'b0101000000001001;    // h364_3=(0.62527)
          9'b101101100:  DATA = 16'b0100111110010010;    // h365_3=(0.62164)
          9'b101101101:  DATA = 16'b0100111100011100;    // h366_3=(0.61804)
          9'b101101110:  DATA = 16'b0100111010100101;    // h367_3=(0.61441)
          9'b101101111:  DATA = 16'b0100111000101101;    // h368_3=(0.61075)
          9'b101110000:  DATA = 16'b0100110110110110;    // h369_3=(0.60712)
          9'b101110001:  DATA = 16'b0100110100111111;    // h370_3=(0.60349)
          9'b101110010:  DATA = 16'b0100110011000111;    // h371_3=(0.59982)
          9'b101110011:  DATA = 16'b0100110001001111;    // h372_3=(0.59616)
          9'b101110100:  DATA = 16'b0100101111010111;    // h373_3=(0.5925)
          9'b101110101:  DATA = 16'b0100101101011111;    // h374_3=(0.58884)
          9'b101110110:  DATA = 16'b0100101011100110;    // h375_3=(0.58514)
          default : DATA = 16'b0000000000000000;
        endcase
    end
endmodule

