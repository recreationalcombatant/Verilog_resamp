`timescale 1ns / 1ps
///////////////////////////////////////////
// ROM table - 2's complement coefficients
// fir_rom4.v: FIR polyphase branch (4)
// 
// Created: 03-Aug-2006 17:33:00
//  from Matlab script fpga_create_rom_verilog.m
//
// J. Shima
//////////////////////////////////////////
module fir_rom4(ADDR, DATA);
    input [8:0] ADDR;
    output signed [15:0] DATA;
    reg signed [15:0] DATA;

    always@(ADDR) begin
        case(ADDR)
          9'b000000000:  DATA = 16'b0100101001101110;    // h1_4=(0.58148)
          9'b000000001:  DATA = 16'b0100100111110101;    // h2_4=(0.57779)
          9'b000000010:  DATA = 16'b0100100101111100;    // h3_4=(0.5741)
          9'b000000011:  DATA = 16'b0100100100000100;    // h4_4=(0.57043)
          9'b000000100:  DATA = 16'b0100100010001010;    // h5_4=(0.56671)
          9'b000000101:  DATA = 16'b0100100000010001;    // h6_4=(0.56302)
          9'b000000110:  DATA = 16'b0100011110011000;    // h7_4=(0.55933)
          9'b000000111:  DATA = 16'b0100011100011111;    // h8_4=(0.55563)
          9'b000001000:  DATA = 16'b0100011010100101;    // h9_4=(0.55191)
          9'b000001001:  DATA = 16'b0100011000101100;    // h10_4=(0.54822)
          9'b000001010:  DATA = 16'b0100010110110010;    // h11_4=(0.54449)
          9'b000001011:  DATA = 16'b0100010100111001;    // h12_4=(0.5408)
          9'b000001100:  DATA = 16'b0100010010111111;    // h13_4=(0.53708)
          9'b000001101:  DATA = 16'b0100010001000101;    // h14_4=(0.53336)
          9'b000001110:  DATA = 16'b0100001111001011;    // h15_4=(0.52963)
          9'b000001111:  DATA = 16'b0100001101010001;    // h16_4=(0.52591)
          9'b000010000:  DATA = 16'b0100001011010111;    // h17_4=(0.52219)
          9'b000010001:  DATA = 16'b0100001001011101;    // h18_4=(0.51846)
          9'b000010010:  DATA = 16'b0100000111100011;    // h19_4=(0.51474)
          9'b000010011:  DATA = 16'b0100000101101001;    // h20_4=(0.51102)
          9'b000010100:  DATA = 16'b0100000011101111;    // h21_4=(0.50729)
          9'b000010101:  DATA = 16'b0100000001110101;    // h22_4=(0.50357)
          9'b000010110:  DATA = 16'b0011111111111011;    // h23_4=(0.49985)
          9'b000010111:  DATA = 16'b0011111110000001;    // h24_4=(0.49612)
          9'b000011000:  DATA = 16'b0011111100000111;    // h25_4=(0.4924)
          9'b000011001:  DATA = 16'b0011111010001101;    // h26_4=(0.48868)
          9'b000011010:  DATA = 16'b0011111000010011;    // h27_4=(0.48495)
          9'b000011011:  DATA = 16'b0011110110011001;    // h28_4=(0.48123)
          9'b000011100:  DATA = 16'b0011110100011111;    // h29_4=(0.47751)
          9'b000011101:  DATA = 16'b0011110010100101;    // h30_4=(0.47379)
          9'b000011110:  DATA = 16'b0011110000101011;    // h31_4=(0.47006)
          9'b000011111:  DATA = 16'b0011101110110001;    // h32_4=(0.46634)
          9'b000100000:  DATA = 16'b0011101100111000;    // h33_4=(0.46265)
          9'b000100001:  DATA = 16'b0011101010111110;    // h34_4=(0.45892)
          9'b000100010:  DATA = 16'b0011101001000100;    // h35_4=(0.4552)
          9'b000100011:  DATA = 16'b0011100111001011;    // h36_4=(0.45151)
          9'b000100100:  DATA = 16'b0011100101010001;    // h37_4=(0.44778)
          9'b000100101:  DATA = 16'b0011100011011000;    // h38_4=(0.44409)
          9'b000100110:  DATA = 16'b0011100001011110;    // h39_4=(0.44037)
          9'b000100111:  DATA = 16'b0011011111100101;    // h40_4=(0.43668)
          9'b000101000:  DATA = 16'b0011011101101100;    // h41_4=(0.43298)
          9'b000101001:  DATA = 16'b0011011011110011;    // h42_4=(0.42929)
          9'b000101010:  DATA = 16'b0011011001111010;    // h43_4=(0.4256)
          9'b000101011:  DATA = 16'b0011011000000001;    // h44_4=(0.42191)
          9'b000101100:  DATA = 16'b0011010110001001;    // h45_4=(0.41824)
          9'b000101101:  DATA = 16'b0011010100010000;    // h46_4=(0.41455)
          9'b000101110:  DATA = 16'b0011010010011000;    // h47_4=(0.41089)
          9'b000101111:  DATA = 16'b0011010000011111;    // h48_4=(0.4072)
          9'b000110000:  DATA = 16'b0011001110100111;    // h49_4=(0.40353)
          9'b000110001:  DATA = 16'b0011001100101111;    // h50_4=(0.39987)
          9'b000110010:  DATA = 16'b0011001010111000;    // h51_4=(0.39624)
          9'b000110011:  DATA = 16'b0011001001000000;    // h52_4=(0.39258)
          9'b000110100:  DATA = 16'b0011000111001000;    // h53_4=(0.38892)
          9'b000110101:  DATA = 16'b0011000101010001;    // h54_4=(0.38528)
          9'b000110110:  DATA = 16'b0011000011011010;    // h55_4=(0.38165)
          9'b000110111:  DATA = 16'b0011000001100011;    // h56_4=(0.37802)
          9'b000111000:  DATA = 16'b0010111111101100;    // h57_4=(0.37439)
          9'b000111001:  DATA = 16'b0010111101110110;    // h58_4=(0.37079)
          9'b000111010:  DATA = 16'b0010111100000000;    // h59_4=(0.36719)
          9'b000111011:  DATA = 16'b0010111010001010;    // h60_4=(0.36359)
          9'b000111100:  DATA = 16'b0010111000010100;    // h61_4=(0.35999)
          9'b000111101:  DATA = 16'b0010110110011110;    // h62_4=(0.35638)
          9'b000111110:  DATA = 16'b0010110100101000;    // h63_4=(0.35278)
          9'b000111111:  DATA = 16'b0010110010110011;    // h64_4=(0.34921)
          9'b001000000:  DATA = 16'b0010110000111110;    // h65_4=(0.34564)
          9'b001000001:  DATA = 16'b0010101111001010;    // h66_4=(0.3421)
          9'b001000010:  DATA = 16'b0010101101010101;    // h67_4=(0.33853)
          9'b001000011:  DATA = 16'b0010101011100001;    // h68_4=(0.33499)
          9'b001000100:  DATA = 16'b0010101001101101;    // h69_4=(0.33145)
          9'b001000101:  DATA = 16'b0010100111111001;    // h70_4=(0.32791)
          9'b001000110:  DATA = 16'b0010100110000110;    // h71_4=(0.3244)
          9'b001000111:  DATA = 16'b0010100100010010;    // h72_4=(0.32086)
          9'b001001000:  DATA = 16'b0010100010011111;    // h73_4=(0.31735)
          9'b001001001:  DATA = 16'b0010100000101101;    // h74_4=(0.31387)
          9'b001001010:  DATA = 16'b0010011110111010;    // h75_4=(0.31036)
          9'b001001011:  DATA = 16'b0010011101001000;    // h76_4=(0.30688)
          9'b001001100:  DATA = 16'b0010011011010111;    // h77_4=(0.30344)
          9'b001001101:  DATA = 16'b0010011001100101;    // h78_4=(0.29996)
          9'b001001110:  DATA = 16'b0010010111110100;    // h79_4=(0.29651)
          9'b001001111:  DATA = 16'b0010010110000011;    // h80_4=(0.29306)
          9'b001010000:  DATA = 16'b0010010100010010;    // h81_4=(0.28961)
          9'b001010001:  DATA = 16'b0010010010100010;    // h82_4=(0.28619)
          9'b001010010:  DATA = 16'b0010010000110010;    // h83_4=(0.28278)
          9'b001010011:  DATA = 16'b0010001111000011;    // h84_4=(0.27939)
          9'b001010100:  DATA = 16'b0010001101010011;    // h85_4=(0.27597)
          9'b001010101:  DATA = 16'b0010001011100100;    // h86_4=(0.27258)
          9'b001010110:  DATA = 16'b0010001001110110;    // h87_4=(0.26923)
          9'b001010111:  DATA = 16'b0010001000001000;    // h88_4=(0.26587)
          9'b001011000:  DATA = 16'b0010000110011010;    // h89_4=(0.26251)
          9'b001011001:  DATA = 16'b0010000100101100;    // h90_4=(0.25916)
          9'b001011010:  DATA = 16'b0010000010111111;    // h91_4=(0.25583)
          9'b001011011:  DATA = 16'b0010000001010010;    // h92_4=(0.2525)
          9'b001011100:  DATA = 16'b0001111111100110;    // h93_4=(0.24921)
          9'b001011101:  DATA = 16'b0001111101111010;    // h94_4=(0.24591)
          9'b001011110:  DATA = 16'b0001111100001110;    // h95_4=(0.24261)
          9'b001011111:  DATA = 16'b0001111010100011;    // h96_4=(0.23935)
          9'b001100000:  DATA = 16'b0001111000111000;    // h97_4=(0.23608)
          9'b001100001:  DATA = 16'b0001110111001101;    // h98_4=(0.23282)
          9'b001100010:  DATA = 16'b0001110101100011;    // h99_4=(0.22958)
          9'b001100011:  DATA = 16'b0001110011111001;    // h100_4=(0.22635)
          9'b001100100:  DATA = 16'b0001110010010000;    // h101_4=(0.22314)
          9'b001100101:  DATA = 16'b0001110000100111;    // h102_4=(0.21994)
          9'b001100110:  DATA = 16'b0001101110111110;    // h103_4=(0.21674)
          9'b001100111:  DATA = 16'b0001101101010110;    // h104_4=(0.21356)
          9'b001101000:  DATA = 16'b0001101011101110;    // h105_4=(0.21039)
          9'b001101001:  DATA = 16'b0001101010000111;    // h106_4=(0.20724)
          9'b001101010:  DATA = 16'b0001101000100000;    // h107_4=(0.2041)
          9'b001101011:  DATA = 16'b0001100110111010;    // h108_4=(0.20099)
          9'b001101100:  DATA = 16'b0001100101010100;    // h109_4=(0.19788)
          9'b001101101:  DATA = 16'b0001100011101110;    // h110_4=(0.19476)
          9'b001101110:  DATA = 16'b0001100010001001;    // h111_4=(0.19168)
          9'b001101111:  DATA = 16'b0001100000100100;    // h112_4=(0.1886)
          9'b001110000:  DATA = 16'b0001011111000000;    // h113_4=(0.18555)
          9'b001110001:  DATA = 16'b0001011101011100;    // h114_4=(0.1825)
          9'b001110010:  DATA = 16'b0001011011111000;    // h115_4=(0.17944)
          9'b001110011:  DATA = 16'b0001011010010101;    // h116_4=(0.17642)
          9'b001110100:  DATA = 16'b0001011000110011;    // h117_4=(0.17343)
          9'b001110101:  DATA = 16'b0001010111010001;    // h118_4=(0.17044)
          9'b001110110:  DATA = 16'b0001010101101111;    // h119_4=(0.16745)
          9'b001110111:  DATA = 16'b0001010100001110;    // h120_4=(0.16449)
          9'b001111000:  DATA = 16'b0001010010101101;    // h121_4=(0.16153)
          9'b001111001:  DATA = 16'b0001010001001101;    // h122_4=(0.1586)
          9'b001111010:  DATA = 16'b0001001111101110;    // h123_4=(0.1557)
          9'b001111011:  DATA = 16'b0001001110001110;    // h124_4=(0.15277)
          9'b001111100:  DATA = 16'b0001001100110000;    // h125_4=(0.1499)
          9'b001111101:  DATA = 16'b0001001011010001;    // h126_4=(0.147)
          9'b001111110:  DATA = 16'b0001001001110011;    // h127_4=(0.14413)
          9'b001111111:  DATA = 16'b0001001000010110;    // h128_4=(0.1413)
          9'b010000000:  DATA = 16'b0001000110111001;    // h129_4=(0.13846)
          9'b010000001:  DATA = 16'b0001000101011101;    // h130_4=(0.13565)
          9'b010000010:  DATA = 16'b0001000100000001;    // h131_4=(0.13284)
          9'b010000011:  DATA = 16'b0001000010100110;    // h132_4=(0.13007)
          9'b010000100:  DATA = 16'b0001000001001011;    // h133_4=(0.12729)
          9'b010000101:  DATA = 16'b0000111111110001;    // h134_4=(0.12454)
          9'b010000110:  DATA = 16'b0000111110010111;    // h135_4=(0.1218)
          9'b010000111:  DATA = 16'b0000111100111101;    // h136_4=(0.11905)
          9'b010001000:  DATA = 16'b0000111011100101;    // h137_4=(0.11636)
          9'b010001001:  DATA = 16'b0000111010001100;    // h138_4=(0.11365)
          9'b010001010:  DATA = 16'b0000111000110101;    // h139_4=(0.11099)
          9'b010001011:  DATA = 16'b0000110111011101;    // h140_4=(0.10831)
          9'b010001100:  DATA = 16'b0000110110000110;    // h141_4=(0.10565)
          9'b010001101:  DATA = 16'b0000110100110000;    // h142_4=(0.10303)
          9'b010001110:  DATA = 16'b0000110011011011;    // h143_4=(0.10043)
          9'b010001111:  DATA = 16'b0000110010000101;    // h144_4=(0.097809)
          9'b010010000:  DATA = 16'b0000110000110001;    // h145_4=(0.095245)
          9'b010010001:  DATA = 16'b0000101111011101;    // h146_4=(0.092682)
          9'b010010010:  DATA = 16'b0000101110001001;    // h147_4=(0.090118)
          9'b010010011:  DATA = 16'b0000101100110110;    // h148_4=(0.087585)
          9'b010010100:  DATA = 16'b0000101011100011;    // h149_4=(0.085052)
          9'b010010101:  DATA = 16'b0000101010010001;    // h150_4=(0.08255)
          9'b010010110:  DATA = 16'b0000101001000000;    // h151_4=(0.080078)
          9'b010010111:  DATA = 16'b0000100111101111;    // h152_4=(0.077606)
          9'b010011000:  DATA = 16'b0000100110011111;    // h153_4=(0.075165)
          9'b010011001:  DATA = 16'b0000100101001111;    // h154_4=(0.072723)
          9'b010011010:  DATA = 16'b0000100100000000;    // h155_4=(0.070313)
          9'b010011011:  DATA = 16'b0000100010110001;    // h156_4=(0.067902)
          9'b010011100:  DATA = 16'b0000100001100011;    // h157_4=(0.065521)
          9'b010011101:  DATA = 16'b0000100000010101;    // h158_4=(0.063141)
          9'b010011110:  DATA = 16'b0000011111001000;    // h159_4=(0.060791)
          9'b010011111:  DATA = 16'b0000011101111011;    // h160_4=(0.058441)
          9'b010100000:  DATA = 16'b0000011100101111;    // h161_4=(0.056122)
          9'b010100001:  DATA = 16'b0000011011100100;    // h162_4=(0.053833)
          9'b010100010:  DATA = 16'b0000011010011001;    // h163_4=(0.051544)
          9'b010100011:  DATA = 16'b0000011001001111;    // h164_4=(0.049286)
          9'b010100100:  DATA = 16'b0000011000000101;    // h165_4=(0.047028)
          9'b010100101:  DATA = 16'b0000010110111100;    // h166_4=(0.0448)
          9'b010100110:  DATA = 16'b0000010101110011;    // h167_4=(0.042572)
          9'b010100111:  DATA = 16'b0000010100101011;    // h168_4=(0.040375)
          9'b010101000:  DATA = 16'b0000010011100011;    // h169_4=(0.038177)
          9'b010101001:  DATA = 16'b0000010010011100;    // h170_4=(0.036011)
          9'b010101010:  DATA = 16'b0000010001010110;    // h171_4=(0.033875)
          9'b010101011:  DATA = 16'b0000010000010000;    // h172_4=(0.031738)
          9'b010101100:  DATA = 16'b0000001111001011;    // h173_4=(0.029633)
          9'b010101101:  DATA = 16'b0000001110000110;    // h174_4=(0.027527)
          9'b010101110:  DATA = 16'b0000001101000010;    // h175_4=(0.025452)
          9'b010101111:  DATA = 16'b0000001011111111;    // h176_4=(0.023407)
          9'b010110000:  DATA = 16'b0000001010111100;    // h177_4=(0.021362)
          9'b010110001:  DATA = 16'b0000001001111001;    // h178_4=(0.019318)
          9'b010110010:  DATA = 16'b0000001000110111;    // h179_4=(0.017303)
          9'b010110011:  DATA = 16'b0000000111110110;    // h180_4=(0.01532)
          9'b010110100:  DATA = 16'b0000000110110101;    // h181_4=(0.013336)
          9'b010110101:  DATA = 16'b0000000101110101;    // h182_4=(0.011383)
          9'b010110110:  DATA = 16'b0000000100110101;    // h183_4=(0.0094299)
          9'b010110111:  DATA = 16'b0000000011110110;    // h184_4=(0.0075073)
          9'b010111000:  DATA = 16'b0000000010111000;    // h185_4=(0.0056152)
          9'b010111001:  DATA = 16'b0000000001111010;    // h186_4=(0.0037231)
          9'b010111010:  DATA = 16'b0000000000111101;    // h187_4=(0.0018616)
          9'b010111011:  DATA = 16'b0000000000000000;    // h188_4=(0)
          9'b010111100:  DATA = 16'b1111111111000100;    // h189_4=(-0.0018311)
          9'b010111101:  DATA = 16'b1111111110001000;    // h190_4=(-0.0036621)
          9'b010111110:  DATA = 16'b1111111101001101;    // h191_4=(-0.0054626)
          9'b010111111:  DATA = 16'b1111111100010011;    // h192_4=(-0.0072327)
          9'b011000000:  DATA = 16'b1111111011011001;    // h193_4=(-0.0090027)
          9'b011000001:  DATA = 16'b1111111010100000;    // h194_4=(-0.010742)
          9'b011000010:  DATA = 16'b1111111001100111;    // h195_4=(-0.012482)
          9'b011000011:  DATA = 16'b1111111000101111;    // h196_4=(-0.014191)
          9'b011000100:  DATA = 16'b1111110111110111;    // h197_4=(-0.0159)
          9'b011000101:  DATA = 16'b1111110111000000;    // h198_4=(-0.017578)
          9'b011000110:  DATA = 16'b1111110110001010;    // h199_4=(-0.019226)
          9'b011000111:  DATA = 16'b1111110101010100;    // h200_4=(-0.020874)
          9'b011001000:  DATA = 16'b1111110100011110;    // h201_4=(-0.022522)
          9'b011001001:  DATA = 16'b1111110011101010;    // h202_4=(-0.024109)
          9'b011001010:  DATA = 16'b1111110010110101;    // h203_4=(-0.025726)
          9'b011001011:  DATA = 16'b1111110010000010;    // h204_4=(-0.027283)
          9'b011001100:  DATA = 16'b1111110001001111;    // h205_4=(-0.028839)
          9'b011001101:  DATA = 16'b1111110000011100;    // h206_4=(-0.030396)
          9'b011001110:  DATA = 16'b1111101111101010;    // h207_4=(-0.031921)
          9'b011001111:  DATA = 16'b1111101110111001;    // h208_4=(-0.033417)
          9'b011010000:  DATA = 16'b1111101110001000;    // h209_4=(-0.034912)
          9'b011010001:  DATA = 16'b1111101101011000;    // h210_4=(-0.036377)
          9'b011010010:  DATA = 16'b1111101100101000;    // h211_4=(-0.037842)
          9'b011010011:  DATA = 16'b1111101011111001;    // h212_4=(-0.039276)
          9'b011010100:  DATA = 16'b1111101011001011;    // h213_4=(-0.04068)
          9'b011010101:  DATA = 16'b1111101010011101;    // h214_4=(-0.042084)
          9'b011010110:  DATA = 16'b1111101001101111;    // h215_4=(-0.043488)
          9'b011010111:  DATA = 16'b1111101001000010;    // h216_4=(-0.044861)
          9'b011011000:  DATA = 16'b1111101000010110;    // h217_4=(-0.046204)
          9'b011011001:  DATA = 16'b1111100111101010;    // h218_4=(-0.047546)
          9'b011011010:  DATA = 16'b1111100110111111;    // h219_4=(-0.048859)
          9'b011011011:  DATA = 16'b1111100110010100;    // h220_4=(-0.050171)
          9'b011011100:  DATA = 16'b1111100101101010;    // h221_4=(-0.051453)
          9'b011011101:  DATA = 16'b1111100101000001;    // h222_4=(-0.052704)
          9'b011011110:  DATA = 16'b1111100100011000;    // h223_4=(-0.053955)
          9'b011011111:  DATA = 16'b1111100011101111;    // h224_4=(-0.055206)
          9'b011100000:  DATA = 16'b1111100011001000;    // h225_4=(-0.056396)
          9'b011100001:  DATA = 16'b1111100010100000;    // h226_4=(-0.057617)
          9'b011100010:  DATA = 16'b1111100001111001;    // h227_4=(-0.058807)
          9'b011100011:  DATA = 16'b1111100001010011;    // h228_4=(-0.059967)
          9'b011100100:  DATA = 16'b1111100000101101;    // h229_4=(-0.061127)
          9'b011100101:  DATA = 16'b1111100000001000;    // h230_4=(-0.062256)
          9'b011100110:  DATA = 16'b1111011111100100;    // h231_4=(-0.063354)
          9'b011100111:  DATA = 16'b1111011111000000;    // h232_4=(-0.064453)
          9'b011101000:  DATA = 16'b1111011110011100;    // h233_4=(-0.065552)
          9'b011101001:  DATA = 16'b1111011101111001;    // h234_4=(-0.06662)
          9'b011101010:  DATA = 16'b1111011101010111;    // h235_4=(-0.067657)
          9'b011101011:  DATA = 16'b1111011100110101;    // h236_4=(-0.068695)
          9'b011101100:  DATA = 16'b1111011100010011;    // h237_4=(-0.069733)
          9'b011101101:  DATA = 16'b1111011011110010;    // h238_4=(-0.07074)
          9'b011101110:  DATA = 16'b1111011011010010;    // h239_4=(-0.071716)
          9'b011101111:  DATA = 16'b1111011010110010;    // h240_4=(-0.072693)
          9'b011110000:  DATA = 16'b1111011010010011;    // h241_4=(-0.073639)
          9'b011110001:  DATA = 16'b1111011001110100;    // h242_4=(-0.074585)
          9'b011110010:  DATA = 16'b1111011001010110;    // h243_4=(-0.0755)
          9'b011110011:  DATA = 16'b1111011000111000;    // h244_4=(-0.076416)
          9'b011110100:  DATA = 16'b1111011000011011;    // h245_4=(-0.077301)
          9'b011110101:  DATA = 16'b1111010111111110;    // h246_4=(-0.078186)
          9'b011110110:  DATA = 16'b1111010111100010;    // h247_4=(-0.079041)
          9'b011110111:  DATA = 16'b1111010111000110;    // h248_4=(-0.079895)
          9'b011111000:  DATA = 16'b1111010110101011;    // h249_4=(-0.080719)
          9'b011111001:  DATA = 16'b1111010110010000;    // h250_4=(-0.081543)
          9'b011111010:  DATA = 16'b1111010101110110;    // h251_4=(-0.082336)
          9'b011111011:  DATA = 16'b1111010101011100;    // h252_4=(-0.08313)
          9'b011111100:  DATA = 16'b1111010101000011;    // h253_4=(-0.083893)
          9'b011111101:  DATA = 16'b1111010100101011;    // h254_4=(-0.084625)
          9'b011111110:  DATA = 16'b1111010100010010;    // h255_4=(-0.085388)
          9'b011111111:  DATA = 16'b1111010011111011;    // h256_4=(-0.08609)
          9'b100000000:  DATA = 16'b1111010011100011;    // h257_4=(-0.086823)
          9'b100000001:  DATA = 16'b1111010011001101;    // h258_4=(-0.087494)
          9'b100000010:  DATA = 16'b1111010010110111;    // h259_4=(-0.088165)
          9'b100000011:  DATA = 16'b1111010010100001;    // h260_4=(-0.088837)
          9'b100000100:  DATA = 16'b1111010010001100;    // h261_4=(-0.089478)
          9'b100000101:  DATA = 16'b1111010001110111;    // h262_4=(-0.090118)
          9'b100000110:  DATA = 16'b1111010001100010;    // h263_4=(-0.090759)
          9'b100000111:  DATA = 16'b1111010001001111;    // h264_4=(-0.091339)
          9'b100001000:  DATA = 16'b1111010000111011;    // h265_4=(-0.091949)
          9'b100001001:  DATA = 16'b1111010000101000;    // h266_4=(-0.092529)
          9'b100001010:  DATA = 16'b1111010000010110;    // h267_4=(-0.093079)
          9'b100001011:  DATA = 16'b1111010000000100;    // h268_4=(-0.093628)
          9'b100001100:  DATA = 16'b1111001111110011;    // h269_4=(-0.094147)
          9'b100001101:  DATA = 16'b1111001111100010;    // h270_4=(-0.094666)
          9'b100001110:  DATA = 16'b1111001111010001;    // h271_4=(-0.095184)
          9'b100001111:  DATA = 16'b1111001111000001;    // h272_4=(-0.095673)
          9'b100010000:  DATA = 16'b1111001110110001;    // h273_4=(-0.096161)
          9'b100010001:  DATA = 16'b1111001110100010;    // h274_4=(-0.096619)
          9'b100010010:  DATA = 16'b1111001110010011;    // h275_4=(-0.097076)
          9'b100010011:  DATA = 16'b1111001110000101;    // h276_4=(-0.097504)
          9'b100010100:  DATA = 16'b1111001101110111;    // h277_4=(-0.097931)
          9'b100010101:  DATA = 16'b1111001101101010;    // h278_4=(-0.098328)
          9'b100010110:  DATA = 16'b1111001101011101;    // h279_4=(-0.098724)
          9'b100010111:  DATA = 16'b1111001101010000;    // h280_4=(-0.099121)
          9'b100011000:  DATA = 16'b1111001101000100;    // h281_4=(-0.099487)
          9'b100011001:  DATA = 16'b1111001100111000;    // h282_4=(-0.099854)
          9'b100011010:  DATA = 16'b1111001100101101;    // h283_4=(-0.10019)
          9'b100011011:  DATA = 16'b1111001100100010;    // h284_4=(-0.10052)
          9'b100011100:  DATA = 16'b1111001100011000;    // h285_4=(-0.10083)
          9'b100011101:  DATA = 16'b1111001100001110;    // h286_4=(-0.10114)
          9'b100011110:  DATA = 16'b1111001100000100;    // h287_4=(-0.10144)
          9'b100011111:  DATA = 16'b1111001011111011;    // h288_4=(-0.10172)
          9'b100100000:  DATA = 16'b1111001011110010;    // h289_4=(-0.10199)
          9'b100100001:  DATA = 16'b1111001011101010;    // h290_4=(-0.10223)
          9'b100100010:  DATA = 16'b1111001011100010;    // h291_4=(-0.10248)
          9'b100100011:  DATA = 16'b1111001011011010;    // h292_4=(-0.10272)
          9'b100100100:  DATA = 16'b1111001011010011;    // h293_4=(-0.10294)
          9'b100100101:  DATA = 16'b1111001011001100;    // h294_4=(-0.10315)
          9'b100100110:  DATA = 16'b1111001011000110;    // h295_4=(-0.10333)
          9'b100100111:  DATA = 16'b1111001011000000;    // h296_4=(-0.10352)
          9'b100101000:  DATA = 16'b1111001010111010;    // h297_4=(-0.1037)
          9'b100101001:  DATA = 16'b1111001010110101;    // h298_4=(-0.10385)
          9'b100101010:  DATA = 16'b1111001010110000;    // h299_4=(-0.104)
          9'b100101011:  DATA = 16'b1111001010101100;    // h300_4=(-0.10413)
          9'b100101100:  DATA = 16'b1111001010101000;    // h301_4=(-0.10425)
          9'b100101101:  DATA = 16'b1111001010100100;    // h302_4=(-0.10437)
          9'b100101110:  DATA = 16'b1111001010100001;    // h303_4=(-0.10446)
          9'b100101111:  DATA = 16'b1111001010011110;    // h304_4=(-0.10455)
          9'b100110000:  DATA = 16'b1111001010011011;    // h305_4=(-0.10464)
          9'b100110001:  DATA = 16'b1111001010011001;    // h306_4=(-0.10471)
          9'b100110010:  DATA = 16'b1111001010010111;    // h307_4=(-0.10477)
          9'b100110011:  DATA = 16'b1111001010010101;    // h308_4=(-0.10483)
          9'b100110100:  DATA = 16'b1111001010010100;    // h309_4=(-0.10486)
          9'b100110101:  DATA = 16'b1111001010010011;    // h310_4=(-0.10489)
          9'b100110110:  DATA = 16'b1111001010010011;    // h311_4=(-0.10489)
          9'b100110111:  DATA = 16'b1111001010010011;    // h312_4=(-0.10489)
          9'b100111000:  DATA = 16'b1111001010010011;    // h313_4=(-0.10489)
          9'b100111001:  DATA = 16'b1111001010010011;    // h314_4=(-0.10489)
          9'b100111010:  DATA = 16'b1111001010010100;    // h315_4=(-0.10486)
          9'b100111011:  DATA = 16'b1111001010010101;    // h316_4=(-0.10483)
          9'b100111100:  DATA = 16'b1111001010010111;    // h317_4=(-0.10477)
          9'b100111101:  DATA = 16'b1111001010011001;    // h318_4=(-0.10471)
          9'b100111110:  DATA = 16'b1111001010011011;    // h319_4=(-0.10464)
          9'b100111111:  DATA = 16'b1111001010011101;    // h320_4=(-0.10458)
          9'b101000000:  DATA = 16'b1111001010100000;    // h321_4=(-0.10449)
          9'b101000001:  DATA = 16'b1111001010100011;    // h322_4=(-0.1044)
          9'b101000010:  DATA = 16'b1111001010100110;    // h323_4=(-0.10431)
          9'b101000011:  DATA = 16'b1111001010101010;    // h324_4=(-0.10419)
          9'b101000100:  DATA = 16'b1111001010101110;    // h325_4=(-0.10406)
          9'b101000101:  DATA = 16'b1111001010110010;    // h326_4=(-0.10394)
          9'b101000110:  DATA = 16'b1111001010110111;    // h327_4=(-0.10379)
          9'b101000111:  DATA = 16'b1111001010111100;    // h328_4=(-0.10364)
          9'b101001000:  DATA = 16'b1111001011000001;    // h329_4=(-0.10349)
          9'b101001001:  DATA = 16'b1111001011000110;    // h330_4=(-0.10333)
          9'b101001010:  DATA = 16'b1111001011001100;    // h331_4=(-0.10315)
          9'b101001011:  DATA = 16'b1111001011010010;    // h332_4=(-0.10297)
          9'b101001100:  DATA = 16'b1111001011011000;    // h333_4=(-0.10278)
          9'b101001101:  DATA = 16'b1111001011011111;    // h334_4=(-0.10257)
          9'b101001110:  DATA = 16'b1111001011100110;    // h335_4=(-0.10236)
          9'b101001111:  DATA = 16'b1111001011101101;    // h336_4=(-0.10214)
          9'b101010000:  DATA = 16'b1111001011110100;    // h337_4=(-0.10193)
          9'b101010001:  DATA = 16'b1111001011111100;    // h338_4=(-0.10168)
          9'b101010010:  DATA = 16'b1111001100000100;    // h339_4=(-0.10144)
          9'b101010011:  DATA = 16'b1111001100001100;    // h340_4=(-0.1012)
          9'b101010100:  DATA = 16'b1111001100010100;    // h341_4=(-0.10095)
          9'b101010101:  DATA = 16'b1111001100011101;    // h342_4=(-0.10068)
          9'b101010110:  DATA = 16'b1111001100100101;    // h343_4=(-0.10043)
          9'b101010111:  DATA = 16'b1111001100101111;    // h344_4=(-0.10013)
          9'b101011000:  DATA = 16'b1111001100111000;    // h345_4=(-0.099854)
          9'b101011001:  DATA = 16'b1111001101000001;    // h346_4=(-0.099579)
          9'b101011010:  DATA = 16'b1111001101001011;    // h347_4=(-0.099274)
          9'b101011011:  DATA = 16'b1111001101010101;    // h348_4=(-0.098969)
          9'b101011100:  DATA = 16'b1111001101011111;    // h349_4=(-0.098663)
          9'b101011101:  DATA = 16'b1111001101101010;    // h350_4=(-0.098328)
          9'b101011110:  DATA = 16'b1111001101110101;    // h351_4=(-0.097992)
          9'b101011111:  DATA = 16'b1111001110000000;    // h352_4=(-0.097656)
          9'b101100000:  DATA = 16'b1111001110001011;    // h353_4=(-0.097321)
          9'b101100001:  DATA = 16'b1111001110010110;    // h354_4=(-0.096985)
          9'b101100010:  DATA = 16'b1111001110100001;    // h355_4=(-0.096649)
          9'b101100011:  DATA = 16'b1111001110101101;    // h356_4=(-0.096283)
          9'b101100100:  DATA = 16'b1111001110111001;    // h357_4=(-0.095917)
          9'b101100101:  DATA = 16'b1111001111000101;    // h358_4=(-0.095551)
          9'b101100110:  DATA = 16'b1111001111010010;    // h359_4=(-0.095154)
          9'b101100111:  DATA = 16'b1111001111011110;    // h360_4=(-0.094788)
          9'b101101000:  DATA = 16'b1111001111101011;    // h361_4=(-0.094391)
          9'b101101001:  DATA = 16'b1111001111111000;    // h362_4=(-0.093994)
          9'b101101010:  DATA = 16'b1111010000000101;    // h363_4=(-0.093597)
          9'b101101011:  DATA = 16'b1111010000010010;    // h364_4=(-0.093201)
          9'b101101100:  DATA = 16'b1111010000011111;    // h365_4=(-0.092804)
          9'b101101101:  DATA = 16'b1111010000101101;    // h366_4=(-0.092377)
          9'b101101110:  DATA = 16'b1111010000111011;    // h367_4=(-0.091949)
          9'b101101111:  DATA = 16'b1111010001001001;    // h368_4=(-0.091522)
          9'b101110000:  DATA = 16'b1111010001010111;    // h369_4=(-0.091095)
          9'b101110001:  DATA = 16'b1111010001100101;    // h370_4=(-0.090668)
          9'b101110010:  DATA = 16'b1111010001110011;    // h371_4=(-0.09024)
          9'b101110011:  DATA = 16'b1111010010000010;    // h372_4=(-0.089783)
          9'b101110100:  DATA = 16'b1111010010010001;    // h373_4=(-0.089325)
          9'b101110101:  DATA = 16'b1111010010011111;    // h374_4=(-0.088898)
          9'b101110110:  DATA = 16'b1111010010101110;    // h375_4=(-0.08844)
          default : DATA = 16'b0000000000000000;
        endcase
    end
endmodule

