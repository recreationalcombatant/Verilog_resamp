`timescale 1ns / 1ps
///////////////////////////////////////////
// ROM table - 2's complement coefficients
// fir_rom1.v: FIR polyphase branch (1)
// 
// Created: 03-Aug-2006 17:32:59
//  from Matlab script fpga_create_rom_verilog.m
//
// J. Shima
//////////////////////////////////////////
module fir_rom1(ADDR, DATA);
    input [8:0] ADDR;
    output signed [15:0] DATA;
    reg signed [15:0] DATA;

    always@(ADDR) begin
        case(ADDR)
          9'b000000000:  DATA = 16'b0000000010011010;    // h1_1=(0.0046997)
          9'b000000001:  DATA = 16'b0000000010011100;    // h2_1=(0.0047607)
          9'b000000010:  DATA = 16'b0000000010011110;    // h3_1=(0.0048218)
          9'b000000011:  DATA = 16'b0000000010100000;    // h4_1=(0.0048828)
          9'b000000100:  DATA = 16'b0000000010100011;    // h5_1=(0.0049744)
          9'b000000101:  DATA = 16'b0000000010100101;    // h6_1=(0.0050354)
          9'b000000110:  DATA = 16'b0000000010100111;    // h7_1=(0.0050964)
          9'b000000111:  DATA = 16'b0000000010101001;    // h8_1=(0.0051575)
          9'b000001000:  DATA = 16'b0000000010101011;    // h9_1=(0.0052185)
          9'b000001001:  DATA = 16'b0000000010101110;    // h10_1=(0.0053101)
          9'b000001010:  DATA = 16'b0000000010110000;    // h11_1=(0.0053711)
          9'b000001011:  DATA = 16'b0000000010110010;    // h12_1=(0.0054321)
          9'b000001100:  DATA = 16'b0000000010110100;    // h13_1=(0.0054932)
          9'b000001101:  DATA = 16'b0000000010110111;    // h14_1=(0.0055847)
          9'b000001110:  DATA = 16'b0000000010111001;    // h15_1=(0.0056458)
          9'b000001111:  DATA = 16'b0000000010111011;    // h16_1=(0.0057068)
          9'b000010000:  DATA = 16'b0000000010111101;    // h17_1=(0.0057678)
          9'b000010001:  DATA = 16'b0000000011000000;    // h18_1=(0.0058594)
          9'b000010010:  DATA = 16'b0000000011000010;    // h19_1=(0.0059204)
          9'b000010011:  DATA = 16'b0000000011000100;    // h20_1=(0.0059814)
          9'b000010100:  DATA = 16'b0000000011000110;    // h21_1=(0.0060425)
          9'b000010101:  DATA = 16'b0000000011001001;    // h22_1=(0.006134)
          9'b000010110:  DATA = 16'b0000000011001011;    // h23_1=(0.0061951)
          9'b000010111:  DATA = 16'b0000000011001101;    // h24_1=(0.0062561)
          9'b000011000:  DATA = 16'b0000000011001111;    // h25_1=(0.0063171)
          9'b000011001:  DATA = 16'b0000000011010001;    // h26_1=(0.0063782)
          9'b000011010:  DATA = 16'b0000000011010100;    // h27_1=(0.0064697)
          9'b000011011:  DATA = 16'b0000000011010110;    // h28_1=(0.0065308)
          9'b000011100:  DATA = 16'b0000000011011000;    // h29_1=(0.0065918)
          9'b000011101:  DATA = 16'b0000000011011010;    // h30_1=(0.0066528)
          9'b000011110:  DATA = 16'b0000000011011100;    // h31_1=(0.0067139)
          9'b000011111:  DATA = 16'b0000000011011110;    // h32_1=(0.0067749)
          9'b000100000:  DATA = 16'b0000000011100001;    // h33_1=(0.0068665)
          9'b000100001:  DATA = 16'b0000000011100011;    // h34_1=(0.0069275)
          9'b000100010:  DATA = 16'b0000000011100101;    // h35_1=(0.0069885)
          9'b000100011:  DATA = 16'b0000000011100111;    // h36_1=(0.0070496)
          9'b000100100:  DATA = 16'b0000000011101001;    // h37_1=(0.0071106)
          9'b000100101:  DATA = 16'b0000000011101011;    // h38_1=(0.0071716)
          9'b000100110:  DATA = 16'b0000000011101101;    // h39_1=(0.0072327)
          9'b000100111:  DATA = 16'b0000000011101111;    // h40_1=(0.0072937)
          9'b000101000:  DATA = 16'b0000000011110001;    // h41_1=(0.0073547)
          9'b000101001:  DATA = 16'b0000000011110011;    // h42_1=(0.0074158)
          9'b000101010:  DATA = 16'b0000000011110101;    // h43_1=(0.0074768)
          9'b000101011:  DATA = 16'b0000000011110111;    // h44_1=(0.0075378)
          9'b000101100:  DATA = 16'b0000000011111001;    // h45_1=(0.0075989)
          9'b000101101:  DATA = 16'b0000000011111011;    // h46_1=(0.0076599)
          9'b000101110:  DATA = 16'b0000000011111101;    // h47_1=(0.0077209)
          9'b000101111:  DATA = 16'b0000000011111111;    // h48_1=(0.007782)
          9'b000110000:  DATA = 16'b0000000100000001;    // h49_1=(0.007843)
          9'b000110001:  DATA = 16'b0000000100000011;    // h50_1=(0.0079041)
          9'b000110010:  DATA = 16'b0000000100000101;    // h51_1=(0.0079651)
          9'b000110011:  DATA = 16'b0000000100000111;    // h52_1=(0.0080261)
          9'b000110100:  DATA = 16'b0000000100001001;    // h53_1=(0.0080872)
          9'b000110101:  DATA = 16'b0000000100001010;    // h54_1=(0.0081177)
          9'b000110110:  DATA = 16'b0000000100001100;    // h55_1=(0.0081787)
          9'b000110111:  DATA = 16'b0000000100001110;    // h56_1=(0.0082397)
          9'b000111000:  DATA = 16'b0000000100010000;    // h57_1=(0.0083008)
          9'b000111001:  DATA = 16'b0000000100010001;    // h58_1=(0.0083313)
          9'b000111010:  DATA = 16'b0000000100010011;    // h59_1=(0.0083923)
          9'b000111011:  DATA = 16'b0000000100010101;    // h60_1=(0.0084534)
          9'b000111100:  DATA = 16'b0000000100010110;    // h61_1=(0.0084839)
          9'b000111101:  DATA = 16'b0000000100011000;    // h62_1=(0.0085449)
          9'b000111110:  DATA = 16'b0000000100011001;    // h63_1=(0.0085754)
          9'b000111111:  DATA = 16'b0000000100011011;    // h64_1=(0.0086365)
          9'b001000000:  DATA = 16'b0000000100011100;    // h65_1=(0.008667)
          9'b001000001:  DATA = 16'b0000000100011110;    // h66_1=(0.008728)
          9'b001000010:  DATA = 16'b0000000100011111;    // h67_1=(0.0087585)
          9'b001000011:  DATA = 16'b0000000100100001;    // h68_1=(0.0088196)
          9'b001000100:  DATA = 16'b0000000100100010;    // h69_1=(0.0088501)
          9'b001000101:  DATA = 16'b0000000100100011;    // h70_1=(0.0088806)
          9'b001000110:  DATA = 16'b0000000100100101;    // h71_1=(0.0089417)
          9'b001000111:  DATA = 16'b0000000100100110;    // h72_1=(0.0089722)
          9'b001001000:  DATA = 16'b0000000100100111;    // h73_1=(0.0090027)
          9'b001001001:  DATA = 16'b0000000100101000;    // h74_1=(0.0090332)
          9'b001001010:  DATA = 16'b0000000100101010;    // h75_1=(0.0090942)
          9'b001001011:  DATA = 16'b0000000100101011;    // h76_1=(0.0091248)
          9'b001001100:  DATA = 16'b0000000100101100;    // h77_1=(0.0091553)
          9'b001001101:  DATA = 16'b0000000100101101;    // h78_1=(0.0091858)
          9'b001001110:  DATA = 16'b0000000100101110;    // h79_1=(0.0092163)
          9'b001001111:  DATA = 16'b0000000100101111;    // h80_1=(0.0092468)
          9'b001010000:  DATA = 16'b0000000100110000;    // h81_1=(0.0092773)
          9'b001010001:  DATA = 16'b0000000100110001;    // h82_1=(0.0093079)
          9'b001010010:  DATA = 16'b0000000100110001;    // h83_1=(0.0093079)
          9'b001010011:  DATA = 16'b0000000100110010;    // h84_1=(0.0093384)
          9'b001010100:  DATA = 16'b0000000100110011;    // h85_1=(0.0093689)
          9'b001010101:  DATA = 16'b0000000100110100;    // h86_1=(0.0093994)
          9'b001010110:  DATA = 16'b0000000100110100;    // h87_1=(0.0093994)
          9'b001010111:  DATA = 16'b0000000100110101;    // h88_1=(0.0094299)
          9'b001011000:  DATA = 16'b0000000100110101;    // h89_1=(0.0094299)
          9'b001011001:  DATA = 16'b0000000100110110;    // h90_1=(0.0094604)
          9'b001011010:  DATA = 16'b0000000100110110;    // h91_1=(0.0094604)
          9'b001011011:  DATA = 16'b0000000100110111;    // h92_1=(0.009491)
          9'b001011100:  DATA = 16'b0000000100110111;    // h93_1=(0.009491)
          9'b001011101:  DATA = 16'b0000000100110111;    // h94_1=(0.009491)
          9'b001011110:  DATA = 16'b0000000100111000;    // h95_1=(0.0095215)
          9'b001011111:  DATA = 16'b0000000100111000;    // h96_1=(0.0095215)
          9'b001100000:  DATA = 16'b0000000100111000;    // h97_1=(0.0095215)
          9'b001100001:  DATA = 16'b0000000100111000;    // h98_1=(0.0095215)
          9'b001100010:  DATA = 16'b0000000100111000;    // h99_1=(0.0095215)
          9'b001100011:  DATA = 16'b0000000100111000;    // h100_1=(0.0095215)
          9'b001100100:  DATA = 16'b0000000100111000;    // h101_1=(0.0095215)
          9'b001100101:  DATA = 16'b0000000100111000;    // h102_1=(0.0095215)
          9'b001100110:  DATA = 16'b0000000100111000;    // h103_1=(0.0095215)
          9'b001100111:  DATA = 16'b0000000100110111;    // h104_1=(0.009491)
          9'b001101000:  DATA = 16'b0000000100110111;    // h105_1=(0.009491)
          9'b001101001:  DATA = 16'b0000000100110111;    // h106_1=(0.009491)
          9'b001101010:  DATA = 16'b0000000100110110;    // h107_1=(0.0094604)
          9'b001101011:  DATA = 16'b0000000100110110;    // h108_1=(0.0094604)
          9'b001101100:  DATA = 16'b0000000100110101;    // h109_1=(0.0094299)
          9'b001101101:  DATA = 16'b0000000100110100;    // h110_1=(0.0093994)
          9'b001101110:  DATA = 16'b0000000100110100;    // h111_1=(0.0093994)
          9'b001101111:  DATA = 16'b0000000100110011;    // h112_1=(0.0093689)
          9'b001110000:  DATA = 16'b0000000100110010;    // h113_1=(0.0093384)
          9'b001110001:  DATA = 16'b0000000100110001;    // h114_1=(0.0093079)
          9'b001110010:  DATA = 16'b0000000100110000;    // h115_1=(0.0092773)
          9'b001110011:  DATA = 16'b0000000100101111;    // h116_1=(0.0092468)
          9'b001110100:  DATA = 16'b0000000100101110;    // h117_1=(0.0092163)
          9'b001110101:  DATA = 16'b0000000100101101;    // h118_1=(0.0091858)
          9'b001110110:  DATA = 16'b0000000100101011;    // h119_1=(0.0091248)
          9'b001110111:  DATA = 16'b0000000100101010;    // h120_1=(0.0090942)
          9'b001111000:  DATA = 16'b0000000100101001;    // h121_1=(0.0090637)
          9'b001111001:  DATA = 16'b0000000100100111;    // h122_1=(0.0090027)
          9'b001111010:  DATA = 16'b0000000100100110;    // h123_1=(0.0089722)
          9'b001111011:  DATA = 16'b0000000100100100;    // h124_1=(0.0089111)
          9'b001111100:  DATA = 16'b0000000100100010;    // h125_1=(0.0088501)
          9'b001111101:  DATA = 16'b0000000100100000;    // h126_1=(0.0087891)
          9'b001111110:  DATA = 16'b0000000100011111;    // h127_1=(0.0087585)
          9'b001111111:  DATA = 16'b0000000100011101;    // h128_1=(0.0086975)
          9'b010000000:  DATA = 16'b0000000100011011;    // h129_1=(0.0086365)
          9'b010000001:  DATA = 16'b0000000100011001;    // h130_1=(0.0085754)
          9'b010000010:  DATA = 16'b0000000100010110;    // h131_1=(0.0084839)
          9'b010000011:  DATA = 16'b0000000100010100;    // h132_1=(0.0084229)
          9'b010000100:  DATA = 16'b0000000100010010;    // h133_1=(0.0083618)
          9'b010000101:  DATA = 16'b0000000100001111;    // h134_1=(0.0082703)
          9'b010000110:  DATA = 16'b0000000100001101;    // h135_1=(0.0082092)
          9'b010000111:  DATA = 16'b0000000100001010;    // h136_1=(0.0081177)
          9'b010001000:  DATA = 16'b0000000100001000;    // h137_1=(0.0080566)
          9'b010001001:  DATA = 16'b0000000100000101;    // h138_1=(0.0079651)
          9'b010001010:  DATA = 16'b0000000100000010;    // h139_1=(0.0078735)
          9'b010001011:  DATA = 16'b0000000011111111;    // h140_1=(0.007782)
          9'b010001100:  DATA = 16'b0000000011111100;    // h141_1=(0.0076904)
          9'b010001101:  DATA = 16'b0000000011111001;    // h142_1=(0.0075989)
          9'b010001110:  DATA = 16'b0000000011110110;    // h143_1=(0.0075073)
          9'b010001111:  DATA = 16'b0000000011110010;    // h144_1=(0.0073853)
          9'b010010000:  DATA = 16'b0000000011101111;    // h145_1=(0.0072937)
          9'b010010001:  DATA = 16'b0000000011101011;    // h146_1=(0.0071716)
          9'b010010010:  DATA = 16'b0000000011101000;    // h147_1=(0.0070801)
          9'b010010011:  DATA = 16'b0000000011100100;    // h148_1=(0.006958)
          9'b010010100:  DATA = 16'b0000000011100000;    // h149_1=(0.0068359)
          9'b010010101:  DATA = 16'b0000000011011101;    // h150_1=(0.0067444)
          9'b010010110:  DATA = 16'b0000000011011001;    // h151_1=(0.0066223)
          9'b010010111:  DATA = 16'b0000000011010101;    // h152_1=(0.0065002)
          9'b010011000:  DATA = 16'b0000000011010001;    // h153_1=(0.0063782)
          9'b010011001:  DATA = 16'b0000000011001100;    // h154_1=(0.0062256)
          9'b010011010:  DATA = 16'b0000000011001000;    // h155_1=(0.0061035)
          9'b010011011:  DATA = 16'b0000000011000100;    // h156_1=(0.0059814)
          9'b010011100:  DATA = 16'b0000000010111111;    // h157_1=(0.0058289)
          9'b010011101:  DATA = 16'b0000000010111010;    // h158_1=(0.0056763)
          9'b010011110:  DATA = 16'b0000000010110110;    // h159_1=(0.0055542)
          9'b010011111:  DATA = 16'b0000000010110001;    // h160_1=(0.0054016)
          9'b010100000:  DATA = 16'b0000000010101100;    // h161_1=(0.005249)
          9'b010100001:  DATA = 16'b0000000010100111;    // h162_1=(0.0050964)
          9'b010100010:  DATA = 16'b0000000010100010;    // h163_1=(0.0049438)
          9'b010100011:  DATA = 16'b0000000010011101;    // h164_1=(0.0047913)
          9'b010100100:  DATA = 16'b0000000010010111;    // h165_1=(0.0046082)
          9'b010100101:  DATA = 16'b0000000010010010;    // h166_1=(0.0044556)
          9'b010100110:  DATA = 16'b0000000010001100;    // h167_1=(0.0042725)
          9'b010100111:  DATA = 16'b0000000010000111;    // h168_1=(0.0041199)
          9'b010101000:  DATA = 16'b0000000010000001;    // h169_1=(0.0039368)
          9'b010101001:  DATA = 16'b0000000001111011;    // h170_1=(0.0037537)
          9'b010101010:  DATA = 16'b0000000001110101;    // h171_1=(0.0035706)
          9'b010101011:  DATA = 16'b0000000001101111;    // h172_1=(0.0033875)
          9'b010101100:  DATA = 16'b0000000001101001;    // h173_1=(0.0032043)
          9'b010101101:  DATA = 16'b0000000001100011;    // h174_1=(0.0030212)
          9'b010101110:  DATA = 16'b0000000001011101;    // h175_1=(0.0028381)
          9'b010101111:  DATA = 16'b0000000001010110;    // h176_1=(0.0026245)
          9'b010110000:  DATA = 16'b0000000001001111;    // h177_1=(0.0024109)
          9'b010110001:  DATA = 16'b0000000001001001;    // h178_1=(0.0022278)
          9'b010110010:  DATA = 16'b0000000001000010;    // h179_1=(0.0020142)
          9'b010110011:  DATA = 16'b0000000000111011;    // h180_1=(0.0018005)
          9'b010110100:  DATA = 16'b0000000000110100;    // h181_1=(0.0015869)
          9'b010110101:  DATA = 16'b0000000000101101;    // h182_1=(0.0013733)
          9'b010110110:  DATA = 16'b0000000000100110;    // h183_1=(0.0011597)
          9'b010110111:  DATA = 16'b0000000000011110;    // h184_1=(0.00091553)
          9'b010111000:  DATA = 16'b0000000000010111;    // h185_1=(0.0007019)
          9'b010111001:  DATA = 16'b0000000000001111;    // h186_1=(0.00045776)
          9'b010111010:  DATA = 16'b0000000000001000;    // h187_1=(0.00024414)
          9'b010111011:  DATA = 16'b0000000000000000;    // h188_1=(0)
          9'b010111100:  DATA = 16'b1111111111111000;    // h189_1=(-0.00024414)
          9'b010111101:  DATA = 16'b1111111111110000;    // h190_1=(-0.00048828)
          9'b010111110:  DATA = 16'b1111111111101000;    // h191_1=(-0.00073242)
          9'b010111111:  DATA = 16'b1111111111100000;    // h192_1=(-0.00097656)
          9'b011000000:  DATA = 16'b1111111111010111;    // h193_1=(-0.0012512)
          9'b011000001:  DATA = 16'b1111111111001111;    // h194_1=(-0.0014954)
          9'b011000010:  DATA = 16'b1111111111000110;    // h195_1=(-0.00177)
          9'b011000011:  DATA = 16'b1111111110111110;    // h196_1=(-0.0020142)
          9'b011000100:  DATA = 16'b1111111110110101;    // h197_1=(-0.0022888)
          9'b011000101:  DATA = 16'b1111111110101100;    // h198_1=(-0.0025635)
          9'b011000110:  DATA = 16'b1111111110100011;    // h199_1=(-0.0028381)
          9'b011000111:  DATA = 16'b1111111110011010;    // h200_1=(-0.0031128)
          9'b011001000:  DATA = 16'b1111111110010001;    // h201_1=(-0.0033875)
          9'b011001001:  DATA = 16'b1111111110000111;    // h202_1=(-0.0036926)
          9'b011001010:  DATA = 16'b1111111101111110;    // h203_1=(-0.0039673)
          9'b011001011:  DATA = 16'b1111111101110100;    // h204_1=(-0.0042725)
          9'b011001100:  DATA = 16'b1111111101101011;    // h205_1=(-0.0045471)
          9'b011001101:  DATA = 16'b1111111101100001;    // h206_1=(-0.0048523)
          9'b011001110:  DATA = 16'b1111111101010111;    // h207_1=(-0.0051575)
          9'b011001111:  DATA = 16'b1111111101001101;    // h208_1=(-0.0054626)
          9'b011010000:  DATA = 16'b1111111101000011;    // h209_1=(-0.0057678)
          9'b011010001:  DATA = 16'b1111111100111000;    // h210_1=(-0.0061035)
          9'b011010010:  DATA = 16'b1111111100101110;    // h211_1=(-0.0064087)
          9'b011010011:  DATA = 16'b1111111100100100;    // h212_1=(-0.0067139)
          9'b011010100:  DATA = 16'b1111111100011001;    // h213_1=(-0.0070496)
          9'b011010101:  DATA = 16'b1111111100001110;    // h214_1=(-0.0073853)
          9'b011010110:  DATA = 16'b1111111100000011;    // h215_1=(-0.0077209)
          9'b011010111:  DATA = 16'b1111111011111000;    // h216_1=(-0.0080566)
          9'b011011000:  DATA = 16'b1111111011101101;    // h217_1=(-0.0083923)
          9'b011011001:  DATA = 16'b1111111011100010;    // h218_1=(-0.008728)
          9'b011011010:  DATA = 16'b1111111011010111;    // h219_1=(-0.0090637)
          9'b011011011:  DATA = 16'b1111111011001100;    // h220_1=(-0.0093994)
          9'b011011100:  DATA = 16'b1111111011000000;    // h221_1=(-0.0097656)
          9'b011011101:  DATA = 16'b1111111010110100;    // h222_1=(-0.010132)
          9'b011011110:  DATA = 16'b1111111010101001;    // h223_1=(-0.010468)
          9'b011011111:  DATA = 16'b1111111010011101;    // h224_1=(-0.010834)
          9'b011100000:  DATA = 16'b1111111010010001;    // h225_1=(-0.0112)
          9'b011100001:  DATA = 16'b1111111010000101;    // h226_1=(-0.011566)
          9'b011100010:  DATA = 16'b1111111001111001;    // h227_1=(-0.011932)
          9'b011100011:  DATA = 16'b1111111001101100;    // h228_1=(-0.012329)
          9'b011100100:  DATA = 16'b1111111001100000;    // h229_1=(-0.012695)
          9'b011100101:  DATA = 16'b1111111001010011;    // h230_1=(-0.013092)
          9'b011100110:  DATA = 16'b1111111001000111;    // h231_1=(-0.013458)
          9'b011100111:  DATA = 16'b1111111000111010;    // h232_1=(-0.013855)
          9'b011101000:  DATA = 16'b1111111000101101;    // h233_1=(-0.014252)
          9'b011101001:  DATA = 16'b1111111000100000;    // h234_1=(-0.014648)
          9'b011101010:  DATA = 16'b1111111000010011;    // h235_1=(-0.015045)
          9'b011101011:  DATA = 16'b1111111000000110;    // h236_1=(-0.015442)
          9'b011101100:  DATA = 16'b1111110111111001;    // h237_1=(-0.015839)
          9'b011101101:  DATA = 16'b1111110111101011;    // h238_1=(-0.016266)
          9'b011101110:  DATA = 16'b1111110111011110;    // h239_1=(-0.016663)
          9'b011101111:  DATA = 16'b1111110111010000;    // h240_1=(-0.01709)
          9'b011110000:  DATA = 16'b1111110111000010;    // h241_1=(-0.017517)
          9'b011110001:  DATA = 16'b1111110110110101;    // h242_1=(-0.017914)
          9'b011110010:  DATA = 16'b1111110110100111;    // h243_1=(-0.018341)
          9'b011110011:  DATA = 16'b1111110110011001;    // h244_1=(-0.018768)
          9'b011110100:  DATA = 16'b1111110110001011;    // h245_1=(-0.019196)
          9'b011110101:  DATA = 16'b1111110101111100;    // h246_1=(-0.019653)
          9'b011110110:  DATA = 16'b1111110101101110;    // h247_1=(-0.020081)
          9'b011110111:  DATA = 16'b1111110101100000;    // h248_1=(-0.020508)
          9'b011111000:  DATA = 16'b1111110101010001;    // h249_1=(-0.020966)
          9'b011111001:  DATA = 16'b1111110101000010;    // h250_1=(-0.021423)
          9'b011111010:  DATA = 16'b1111110100110100;    // h251_1=(-0.021851)
          9'b011111011:  DATA = 16'b1111110100100101;    // h252_1=(-0.022308)
          9'b011111100:  DATA = 16'b1111110100010110;    // h253_1=(-0.022766)
          9'b011111101:  DATA = 16'b1111110100000111;    // h254_1=(-0.023224)
          9'b011111110:  DATA = 16'b1111110011111000;    // h255_1=(-0.023682)
          9'b011111111:  DATA = 16'b1111110011101001;    // h256_1=(-0.024139)
          9'b100000000:  DATA = 16'b1111110011011001;    // h257_1=(-0.024628)
          9'b100000001:  DATA = 16'b1111110011001010;    // h258_1=(-0.025085)
          9'b100000010:  DATA = 16'b1111110010111010;    // h259_1=(-0.025574)
          9'b100000011:  DATA = 16'b1111110010101011;    // h260_1=(-0.026031)
          9'b100000100:  DATA = 16'b1111110010011011;    // h261_1=(-0.02652)
          9'b100000101:  DATA = 16'b1111110010001011;    // h262_1=(-0.027008)
          9'b100000110:  DATA = 16'b1111110001111100;    // h263_1=(-0.027466)
          9'b100000111:  DATA = 16'b1111110001101100;    // h264_1=(-0.027954)
          9'b100001000:  DATA = 16'b1111110001011100;    // h265_1=(-0.028442)
          9'b100001001:  DATA = 16'b1111110001001011;    // h266_1=(-0.028961)
          9'b100001010:  DATA = 16'b1111110000111011;    // h267_1=(-0.029449)
          9'b100001011:  DATA = 16'b1111110000101011;    // h268_1=(-0.029938)
          9'b100001100:  DATA = 16'b1111110000011011;    // h269_1=(-0.030426)
          9'b100001101:  DATA = 16'b1111110000001010;    // h270_1=(-0.030945)
          9'b100001110:  DATA = 16'b1111101111111010;    // h271_1=(-0.031433)
          9'b100001111:  DATA = 16'b1111101111101001;    // h272_1=(-0.031952)
          9'b100010000:  DATA = 16'b1111101111011000;    // h273_1=(-0.032471)
          9'b100010001:  DATA = 16'b1111101111000111;    // h274_1=(-0.03299)
          9'b100010010:  DATA = 16'b1111101110110111;    // h275_1=(-0.033478)
          9'b100010011:  DATA = 16'b1111101110100110;    // h276_1=(-0.033997)
          9'b100010100:  DATA = 16'b1111101110010101;    // h277_1=(-0.034515)
          9'b100010101:  DATA = 16'b1111101110000100;    // h278_1=(-0.035034)
          9'b100010110:  DATA = 16'b1111101101110010;    // h279_1=(-0.035583)
          9'b100010111:  DATA = 16'b1111101101100001;    // h280_1=(-0.036102)
          9'b100011000:  DATA = 16'b1111101101010000;    // h281_1=(-0.036621)
          9'b100011001:  DATA = 16'b1111101100111110;    // h282_1=(-0.03717)
          9'b100011010:  DATA = 16'b1111101100101101;    // h283_1=(-0.037689)
          9'b100011011:  DATA = 16'b1111101100011100;    // h284_1=(-0.038208)
          9'b100011100:  DATA = 16'b1111101100001010;    // h285_1=(-0.038757)
          9'b100011101:  DATA = 16'b1111101011111000;    // h286_1=(-0.039307)
          9'b100011110:  DATA = 16'b1111101011100111;    // h287_1=(-0.039825)
          9'b100011111:  DATA = 16'b1111101011010101;    // h288_1=(-0.040375)
          9'b100100000:  DATA = 16'b1111101011000011;    // h289_1=(-0.040924)
          9'b100100001:  DATA = 16'b1111101010110001;    // h290_1=(-0.041473)
          9'b100100010:  DATA = 16'b1111101010011111;    // h291_1=(-0.042023)
          9'b100100011:  DATA = 16'b1111101010001101;    // h292_1=(-0.042572)
          9'b100100100:  DATA = 16'b1111101001111011;    // h293_1=(-0.043121)
          9'b100100101:  DATA = 16'b1111101001101001;    // h294_1=(-0.043671)
          9'b100100110:  DATA = 16'b1111101001010111;    // h295_1=(-0.04422)
          9'b100100111:  DATA = 16'b1111101001000101;    // h296_1=(-0.044769)
          9'b100101000:  DATA = 16'b1111101000110011;    // h297_1=(-0.045319)
          9'b100101001:  DATA = 16'b1111101000100001;    // h298_1=(-0.045868)
          9'b100101010:  DATA = 16'b1111101000001110;    // h299_1=(-0.046448)
          9'b100101011:  DATA = 16'b1111100111111100;    // h300_1=(-0.046997)
          9'b100101100:  DATA = 16'b1111100111101010;    // h301_1=(-0.047546)
          9'b100101101:  DATA = 16'b1111100111010111;    // h302_1=(-0.048126)
          9'b100101110:  DATA = 16'b1111100111000101;    // h303_1=(-0.048676)
          9'b100101111:  DATA = 16'b1111100110110010;    // h304_1=(-0.049255)
          9'b100110000:  DATA = 16'b1111100110100000;    // h305_1=(-0.049805)
          9'b100110001:  DATA = 16'b1111100110001101;    // h306_1=(-0.050385)
          9'b100110010:  DATA = 16'b1111100101111011;    // h307_1=(-0.050934)
          9'b100110011:  DATA = 16'b1111100101101000;    // h308_1=(-0.051514)
          9'b100110100:  DATA = 16'b1111100101010101;    // h309_1=(-0.052094)
          9'b100110101:  DATA = 16'b1111100101000011;    // h310_1=(-0.052643)
          9'b100110110:  DATA = 16'b1111100100110000;    // h311_1=(-0.053223)
          9'b100110111:  DATA = 16'b1111100100011101;    // h312_1=(-0.053802)
          9'b100111000:  DATA = 16'b1111100100001011;    // h313_1=(-0.054352)
          9'b100111001:  DATA = 16'b1111100011111000;    // h314_1=(-0.054932)
          9'b100111010:  DATA = 16'b1111100011100101;    // h315_1=(-0.055511)
          9'b100111011:  DATA = 16'b1111100011010010;    // h316_1=(-0.056091)
          9'b100111100:  DATA = 16'b1111100011000000;    // h317_1=(-0.056641)
          9'b100111101:  DATA = 16'b1111100010101101;    // h318_1=(-0.05722)
          9'b100111110:  DATA = 16'b1111100010011010;    // h319_1=(-0.0578)
          9'b100111111:  DATA = 16'b1111100010000111;    // h320_1=(-0.05838)
          9'b101000000:  DATA = 16'b1111100001110101;    // h321_1=(-0.058929)
          9'b101000001:  DATA = 16'b1111100001100010;    // h322_1=(-0.059509)
          9'b101000010:  DATA = 16'b1111100001001111;    // h323_1=(-0.060089)
          9'b101000011:  DATA = 16'b1111100000111100;    // h324_1=(-0.060669)
          9'b101000100:  DATA = 16'b1111100000101010;    // h325_1=(-0.061218)
          9'b101000101:  DATA = 16'b1111100000010111;    // h326_1=(-0.061798)
          9'b101000110:  DATA = 16'b1111100000000100;    // h327_1=(-0.062378)
          9'b101000111:  DATA = 16'b1111011111110001;    // h328_1=(-0.062958)
          9'b101001000:  DATA = 16'b1111011111011111;    // h329_1=(-0.063507)
          9'b101001001:  DATA = 16'b1111011111001100;    // h330_1=(-0.064087)
          9'b101001010:  DATA = 16'b1111011110111001;    // h331_1=(-0.064667)
          9'b101001011:  DATA = 16'b1111011110100111;    // h332_1=(-0.065216)
          9'b101001100:  DATA = 16'b1111011110010100;    // h333_1=(-0.065796)
          9'b101001101:  DATA = 16'b1111011110000001;    // h334_1=(-0.066376)
          9'b101001110:  DATA = 16'b1111011101101111;    // h335_1=(-0.066925)
          9'b101001111:  DATA = 16'b1111011101011100;    // h336_1=(-0.067505)
          9'b101010000:  DATA = 16'b1111011101001010;    // h337_1=(-0.068054)
          9'b101010001:  DATA = 16'b1111011100110111;    // h338_1=(-0.068634)
          9'b101010010:  DATA = 16'b1111011100100101;    // h339_1=(-0.069183)
          9'b101010011:  DATA = 16'b1111011100010011;    // h340_1=(-0.069733)
          9'b101010100:  DATA = 16'b1111011100000000;    // h341_1=(-0.070313)
          9'b101010101:  DATA = 16'b1111011011101110;    // h342_1=(-0.070862)
          9'b101010110:  DATA = 16'b1111011011011100;    // h343_1=(-0.071411)
          9'b101010111:  DATA = 16'b1111011011001001;    // h344_1=(-0.071991)
          9'b101011000:  DATA = 16'b1111011010110111;    // h345_1=(-0.07254)
          9'b101011001:  DATA = 16'b1111011010100101;    // h346_1=(-0.07309)
          9'b101011010:  DATA = 16'b1111011010010011;    // h347_1=(-0.073639)
          9'b101011011:  DATA = 16'b1111011010000001;    // h348_1=(-0.074188)
          9'b101011100:  DATA = 16'b1111011001101111;    // h349_1=(-0.074738)
          9'b101011101:  DATA = 16'b1111011001011110;    // h350_1=(-0.075256)
          9'b101011110:  DATA = 16'b1111011001001100;    // h351_1=(-0.075806)
          9'b101011111:  DATA = 16'b1111011000111010;    // h352_1=(-0.076355)
          9'b101100000:  DATA = 16'b1111011000101000;    // h353_1=(-0.076904)
          9'b101100001:  DATA = 16'b1111011000010111;    // h354_1=(-0.077423)
          9'b101100010:  DATA = 16'b1111011000000110;    // h355_1=(-0.077942)
          9'b101100011:  DATA = 16'b1111010111110100;    // h356_1=(-0.078491)
          9'b101100100:  DATA = 16'b1111010111100011;    // h357_1=(-0.07901)
          9'b101100101:  DATA = 16'b1111010111010010;    // h358_1=(-0.079529)
          9'b101100110:  DATA = 16'b1111010111000001;    // h359_1=(-0.080048)
          9'b101100111:  DATA = 16'b1111010110110000;    // h360_1=(-0.080566)
          9'b101101000:  DATA = 16'b1111010110011111;    // h361_1=(-0.081085)
          9'b101101001:  DATA = 16'b1111010110001110;    // h362_1=(-0.081604)
          9'b101101010:  DATA = 16'b1111010101111101;    // h363_1=(-0.082123)
          9'b101101011:  DATA = 16'b1111010101101100;    // h364_1=(-0.082642)
          9'b101101100:  DATA = 16'b1111010101011100;    // h365_1=(-0.08313)
          9'b101101101:  DATA = 16'b1111010101001100;    // h366_1=(-0.083618)
          9'b101101110:  DATA = 16'b1111010100111011;    // h367_1=(-0.084137)
          9'b101101111:  DATA = 16'b1111010100101011;    // h368_1=(-0.084625)
          9'b101110000:  DATA = 16'b1111010100011011;    // h369_1=(-0.085114)
          9'b101110001:  DATA = 16'b1111010100001011;    // h370_1=(-0.085602)
          9'b101110010:  DATA = 16'b1111010011111011;    // h371_1=(-0.08609)
          9'b101110011:  DATA = 16'b1111010011101100;    // h372_1=(-0.086548)
          9'b101110100:  DATA = 16'b1111010011011100;    // h373_1=(-0.087036)
          9'b101110101:  DATA = 16'b1111010011001101;    // h374_1=(-0.087494)
          9'b101110110:  DATA = 16'b1111010010111101;    // h375_1=(-0.087982)
          default : DATA = 16'b0000000000000000;
        endcase
    end
endmodule

